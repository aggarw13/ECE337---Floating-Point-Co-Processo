// $Id: $
// File name:   tb_Floating_point_co_processor.sv
// Created:     4/30/2015
// Author:      James Alliger
// Lab Section: 337-05
// Version:     1.0  Initial Design Entry
// Description: The main test bench for the floating point co-processor
