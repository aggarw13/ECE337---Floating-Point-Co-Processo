
module scheduling_logic ( instruction1, dependency, instruction_available, 
        dependency_add, sram_address_store, sram_address_load, source1, 
        source2, read_instruction1, store2_enable, store1_enable, load_enable, 
        add_enable, sub_enable, mul_enable, sin_enable, neg_enable, abs_enable, 
        move_enable, load_dest, add_dest, sub_dest, mul_dest, sin_dest, 
        neg_dest, abs_dest, move_dest );
  input [15:0] instruction1;
  input [15:0] dependency;
  output [15:0] dependency_add;
  output [7:0] sram_address_store;
  output [7:0] sram_address_load;
  output [3:0] source1;
  output [3:0] source2;
  output [3:0] load_dest;
  output [3:0] add_dest;
  output [3:0] sub_dest;
  output [3:0] mul_dest;
  output [3:0] sin_dest;
  output [3:0] neg_dest;
  output [3:0] abs_dest;
  output [3:0] move_dest;
  input instruction_available;
  output read_instruction1, store2_enable, store1_enable, load_enable,
         add_enable, sub_enable, mul_enable, sin_enable, neg_enable,
         abs_enable, move_enable;
  wire   N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n95, n97, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n263, n268, n269, n270, n271, n272;
  assign N50 = instruction1[0];
  assign N51 = instruction1[1];
  assign N52 = instruction1[2];
  assign N53 = instruction1[3];
  assign N54 = instruction1[8];
  assign N55 = instruction1[9];
  assign N56 = instruction1[10];
  assign N57 = instruction1[11];
  assign N58 = instruction1[4];
  assign N59 = instruction1[5];
  assign N60 = instruction1[6];
  assign N61 = instruction1[7];

  AND2X2 U3 ( .A(n141), .B(n198), .Y(n196) );
  AND2X2 U4 ( .A(instruction1[14]), .B(n225), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n200) );
  INVX1 U6 ( .A(n64), .Y(n2) );
  INVX4 U7 ( .A(instruction1[14]), .Y(n202) );
  OR2X2 U8 ( .A(n17), .B(n89), .Y(n11) );
  INVX2 U9 ( .A(N53), .Y(n3) );
  INVX2 U10 ( .A(n3), .Y(n4) );
  INVX2 U11 ( .A(N50), .Y(n217) );
  INVX1 U12 ( .A(n225), .Y(n5) );
  INVX2 U13 ( .A(n237), .Y(n8) );
  BUFX2 U14 ( .A(n73), .Y(n6) );
  INVX1 U15 ( .A(n15), .Y(n7) );
  INVX2 U16 ( .A(n29), .Y(n85) );
  INVX1 U17 ( .A(n219), .Y(n9) );
  INVX1 U18 ( .A(n111), .Y(n10) );
  BUFX4 U19 ( .A(n238), .Y(n17) );
  INVX2 U20 ( .A(n170), .Y(n59) );
  INVX2 U21 ( .A(instruction1[15]), .Y(n225) );
  NAND2X1 U22 ( .A(n12), .B(n13), .Y(n14) );
  NAND2X1 U23 ( .A(n14), .B(n79), .Y(n210) );
  INVX1 U24 ( .A(n42), .Y(n12) );
  INVX2 U25 ( .A(n204), .Y(n13) );
  BUFX2 U26 ( .A(N60), .Y(n15) );
  INVX1 U27 ( .A(n198), .Y(n195) );
  INVX1 U28 ( .A(n252), .Y(n16) );
  INVX1 U29 ( .A(n252), .Y(n255) );
  BUFX2 U30 ( .A(n238), .Y(n84) );
  AND2X2 U31 ( .A(n83), .B(n93), .Y(n18) );
  INVX1 U32 ( .A(n42), .Y(n241) );
  INVX2 U33 ( .A(n141), .Y(n23) );
  INVX1 U34 ( .A(n195), .Y(n19) );
  INVX2 U35 ( .A(n56), .Y(n20) );
  INVX1 U36 ( .A(n191), .Y(n176) );
  AND2X2 U37 ( .A(n168), .B(n21), .Y(n190) );
  NOR2X1 U38 ( .A(n22), .B(n123), .Y(n21) );
  NAND2X1 U39 ( .A(n124), .B(n72), .Y(n22) );
  INVX2 U40 ( .A(n110), .Y(n168) );
  INVX1 U41 ( .A(n39), .Y(n214) );
  AND2X2 U42 ( .A(n23), .B(n170), .Y(n81) );
  INVX1 U43 ( .A(n218), .Y(n24) );
  INVX2 U44 ( .A(N51), .Y(n218) );
  INVX1 U45 ( .A(N57), .Y(n82) );
  AND2X2 U46 ( .A(n54), .B(n31), .Y(n25) );
  AND2X2 U47 ( .A(n93), .B(n54), .Y(n26) );
  INVX2 U48 ( .A(n31), .Y(n93) );
  NAND2X1 U49 ( .A(n34), .B(n25), .Y(n27) );
  INVX1 U50 ( .A(n89), .Y(n28) );
  AND2X2 U51 ( .A(n8), .B(n238), .Y(n29) );
  INVX2 U52 ( .A(N54), .Y(n237) );
  BUFX2 U53 ( .A(N54), .Y(n89) );
  INVX1 U54 ( .A(n87), .Y(n30) );
  INVX1 U55 ( .A(n46), .Y(n260) );
  INVX1 U56 ( .A(n91), .Y(n31) );
  AND2X2 U57 ( .A(instruction1[15]), .B(instruction_available), .Y(n76) );
  NAND2X1 U58 ( .A(n34), .B(n18), .Y(n32) );
  INVX1 U59 ( .A(n2), .Y(n33) );
  NAND2X1 U60 ( .A(n255), .B(n256), .Y(n34) );
  NOR2X1 U61 ( .A(instruction1[13]), .B(instruction1[12]), .Y(n73) );
  INVX1 U62 ( .A(n52), .Y(n186) );
  INVX1 U63 ( .A(instruction1[12]), .Y(n185) );
  INVX1 U64 ( .A(n215), .Y(n201) );
  INVX1 U65 ( .A(n241), .Y(n35) );
  BUFX2 U66 ( .A(n52), .Y(n36) );
  INVX1 U67 ( .A(n9), .Y(n269) );
  INVX2 U68 ( .A(N56), .Y(n91) );
  AND2X2 U69 ( .A(n1), .B(n36), .Y(n37) );
  INVX1 U70 ( .A(n37), .Y(n242) );
  INVX1 U71 ( .A(n249), .Y(mul_enable) );
  BUFX2 U72 ( .A(n81), .Y(n38) );
  NAND2X1 U73 ( .A(n81), .B(n190), .Y(n39) );
  INVX1 U74 ( .A(n65), .Y(n40) );
  BUFX2 U75 ( .A(N57), .Y(n87) );
  INVX4 U76 ( .A(n54), .Y(n83) );
  INVX1 U77 ( .A(n7), .Y(n51) );
  INVX2 U78 ( .A(n175), .Y(n41) );
  OR2X1 U79 ( .A(n213), .B(n214), .Y(read_instruction1) );
  AND2X2 U80 ( .A(n71), .B(n76), .Y(n42) );
  INVX2 U81 ( .A(n28), .Y(n43) );
  INVX1 U82 ( .A(n103), .Y(n44) );
  INVX2 U83 ( .A(N59), .Y(n61) );
  AND2X2 U84 ( .A(n238), .B(n237), .Y(n45) );
  INVX4 U85 ( .A(n45), .Y(n64) );
  INVX2 U86 ( .A(mul_enable), .Y(n95) );
  INVX1 U87 ( .A(n51), .Y(n271) );
  AND2X1 U88 ( .A(n83), .B(n31), .Y(n75) );
  OR2X2 U89 ( .A(n60), .B(N59), .Y(n115) );
  AND2X2 U90 ( .A(N55), .B(N54), .Y(n46) );
  NAND2X1 U91 ( .A(n34), .B(n18), .Y(n253) );
  NAND2X1 U92 ( .A(n34), .B(n25), .Y(n259) );
  NAND2X1 U93 ( .A(n65), .B(n100), .Y(n47) );
  INVX1 U94 ( .A(n44), .Y(n272) );
  INVX1 U95 ( .A(n100), .Y(n48) );
  INVX2 U96 ( .A(N58), .Y(n60) );
  BUFX2 U97 ( .A(n185), .Y(n49) );
  INVX1 U98 ( .A(n40), .Y(n50) );
  INVX2 U99 ( .A(n61), .Y(n65) );
  OR2X2 U100 ( .A(N51), .B(N50), .Y(n161) );
  BUFX4 U101 ( .A(instruction1[13]), .Y(n52) );
  INVX1 U102 ( .A(n48), .Y(n270) );
  NAND2X1 U103 ( .A(n67), .B(n218), .Y(n53) );
  INVX1 U104 ( .A(n30), .Y(n54) );
  INVX2 U105 ( .A(load_enable), .Y(n97) );
  INVX1 U106 ( .A(n245), .Y(load_enable) );
  BUFX2 U107 ( .A(n206), .Y(n55) );
  INVX1 U108 ( .A(n220), .Y(n56) );
  BUFX2 U109 ( .A(n207), .Y(n57) );
  BUFX2 U110 ( .A(n79), .Y(n58) );
  INVX1 U111 ( .A(N58), .Y(n100) );
  OR2X2 U112 ( .A(n84), .B(n8), .Y(n62) );
  OR2X2 U113 ( .A(n17), .B(n89), .Y(n63) );
  BUFX2 U114 ( .A(n86), .Y(n66) );
  INVX1 U115 ( .A(n251), .Y(n175) );
  INVX1 U116 ( .A(n17), .Y(n90) );
  NAND2X1 U117 ( .A(n26), .B(n258), .Y(n257) );
  BUFX2 U118 ( .A(N50), .Y(n67) );
  INVX1 U119 ( .A(n90), .Y(n68) );
  BUFX2 U120 ( .A(n11), .Y(n69) );
  AND2X2 U121 ( .A(N51), .B(N50), .Y(n78) );
  INVX1 U122 ( .A(n193), .Y(n180) );
  AND2X2 U123 ( .A(n142), .B(n37), .Y(n70) );
  AND2X2 U124 ( .A(n73), .B(n202), .Y(n71) );
  AND2X2 U125 ( .A(n76), .B(n202), .Y(n72) );
  AND2X2 U126 ( .A(n175), .B(instruction_available), .Y(n74) );
  AND2X2 U127 ( .A(N59), .B(N58), .Y(n77) );
  AND2X2 U128 ( .A(n167), .B(n168), .Y(n79) );
  AND2X2 U129 ( .A(n23), .B(n170), .Y(n80) );
  INVX2 U130 ( .A(n239), .Y(store2_enable) );
  INVX2 U131 ( .A(n240), .Y(store1_enable) );
  INVX1 U132 ( .A(n24), .Y(n268) );
  INVX1 U133 ( .A(n67), .Y(n263) );
  INVX2 U134 ( .A(N55), .Y(n238) );
  INVX2 U135 ( .A(n29), .Y(n86) );
  BUFX2 U136 ( .A(n66), .Y(n88) );
  NAND2X1 U137 ( .A(n75), .B(n258), .Y(n254) );
  INVX1 U138 ( .A(n31), .Y(n92) );
  NOR2X1 U139 ( .A(n52), .B(n185), .Y(n124) );
  NAND2X1 U140 ( .A(n65), .B(n100), .Y(n114) );
  OAI22X1 U141 ( .A(dependency[5]), .B(n115), .C(dependency[6]), .D(n114), .Y(
        n109) );
  NAND2X1 U142 ( .A(n60), .B(n61), .Y(n118) );
  INVX2 U143 ( .A(dependency[7]), .Y(n154) );
  INVX2 U144 ( .A(N61), .Y(n103) );
  NAND2X1 U145 ( .A(n10), .B(n103), .Y(n101) );
  AOI21X1 U146 ( .A(n154), .B(n77), .C(n101), .Y(n102) );
  OAI21X1 U147 ( .A(dependency[4]), .B(n118), .C(n102), .Y(n108) );
  OAI22X1 U148 ( .A(dependency[1]), .B(n115), .C(dependency[2]), .D(n114), .Y(
        n107) );
  INVX2 U149 ( .A(dependency[3]), .Y(n159) );
  INVX2 U150 ( .A(N60), .Y(n111) );
  NAND2X1 U151 ( .A(n111), .B(n103), .Y(n104) );
  AOI21X1 U152 ( .A(n77), .B(n159), .C(n104), .Y(n105) );
  OAI21X1 U153 ( .A(dependency[0]), .B(n118), .C(n105), .Y(n106) );
  OAI22X1 U154 ( .A(n109), .B(n108), .C(n107), .D(n106), .Y(n110) );
  OAI22X1 U155 ( .A(dependency[9]), .B(n115), .C(dependency[10]), .D(n47), .Y(
        n122) );
  INVX2 U156 ( .A(dependency[11]), .Y(n144) );
  NAND2X1 U157 ( .A(n111), .B(N61), .Y(n112) );
  AOI21X1 U158 ( .A(n77), .B(n144), .C(n112), .Y(n113) );
  OAI21X1 U159 ( .A(dependency[8]), .B(n118), .C(n113), .Y(n121) );
  OAI22X1 U160 ( .A(dependency[13]), .B(n115), .C(dependency[14]), .D(n47), 
        .Y(n120) );
  INVX2 U161 ( .A(dependency[15]), .Y(n147) );
  NAND2X1 U162 ( .A(N61), .B(n15), .Y(n116) );
  AOI21X1 U163 ( .A(n77), .B(n147), .C(n116), .Y(n117) );
  OAI21X1 U164 ( .A(n118), .B(dependency[12]), .C(n117), .Y(n119) );
  OAI22X1 U165 ( .A(n122), .B(n121), .C(n119), .D(n120), .Y(n123) );
  INVX2 U166 ( .A(n123), .Y(n167) );
  OAI22X1 U167 ( .A(dependency[9]), .B(n85), .C(dependency[10]), .D(n62), .Y(
        n132) );
  NAND2X1 U168 ( .A(n87), .B(n91), .Y(n125) );
  AOI21X1 U169 ( .A(n144), .B(n46), .C(n125), .Y(n126) );
  OAI21X1 U170 ( .A(dependency[8]), .B(n64), .C(n126), .Y(n131) );
  OAI22X1 U171 ( .A(dependency[1]), .B(n86), .C(dependency[2]), .D(n11), .Y(
        n130) );
  NAND2X1 U172 ( .A(n82), .B(n91), .Y(n127) );
  AOI21X1 U173 ( .A(n46), .B(n159), .C(n127), .Y(n128) );
  OAI21X1 U174 ( .A(dependency[0]), .B(n64), .C(n128), .Y(n129) );
  OAI22X1 U175 ( .A(n132), .B(n131), .C(n130), .D(n129), .Y(n197) );
  INVX2 U176 ( .A(n197), .Y(n170) );
  OAI22X1 U177 ( .A(dependency[5]), .B(n86), .C(dependency[6]), .D(n62), .Y(
        n140) );
  NAND2X1 U178 ( .A(N56), .B(n82), .Y(n133) );
  AOI21X1 U179 ( .A(n154), .B(n46), .C(n133), .Y(n134) );
  OAI21X1 U180 ( .A(dependency[4]), .B(n64), .C(n134), .Y(n139) );
  OAI22X1 U181 ( .A(dependency[13]), .B(n85), .C(dependency[14]), .D(n63), .Y(
        n138) );
  NAND2X1 U182 ( .A(N56), .B(n87), .Y(n135) );
  AOI21X1 U183 ( .A(n46), .B(n147), .C(n135), .Y(n136) );
  OAI21X1 U184 ( .A(dependency[12]), .B(n64), .C(n136), .Y(n137) );
  OAI22X1 U185 ( .A(n139), .B(n140), .C(n138), .D(n137), .Y(n141) );
  NAND2X1 U186 ( .A(n190), .B(n38), .Y(n227) );
  NOR2X1 U187 ( .A(n28), .B(n227), .Y(move_dest[0]) );
  NOR2X1 U188 ( .A(n68), .B(n227), .Y(move_dest[1]) );
  NOR2X1 U189 ( .A(n92), .B(n227), .Y(move_dest[2]) );
  NOR2X1 U190 ( .A(n83), .B(n227), .Y(move_dest[3]) );
  NAND2X1 U191 ( .A(n38), .B(n58), .Y(n224) );
  INVX2 U192 ( .A(n224), .Y(n142) );
  NAND2X1 U193 ( .A(n35), .B(n142), .Y(n181) );
  NOR2X1 U194 ( .A(n28), .B(n181), .Y(abs_dest[0]) );
  NOR2X1 U195 ( .A(n68), .B(n181), .Y(abs_dest[1]) );
  NOR2X1 U196 ( .A(n92), .B(n181), .Y(abs_dest[2]) );
  NOR2X1 U197 ( .A(n83), .B(n181), .Y(abs_dest[3]) );
  NAND2X1 U198 ( .A(instruction1[12]), .B(instruction_available), .Y(n171) );
  INVX2 U199 ( .A(n171), .Y(n189) );
  NAND2X1 U200 ( .A(n70), .B(n189), .Y(n182) );
  NOR2X1 U201 ( .A(n28), .B(n182), .Y(neg_dest[0]) );
  NOR2X1 U202 ( .A(n68), .B(n182), .Y(neg_dest[1]) );
  NOR2X1 U203 ( .A(n92), .B(n182), .Y(neg_dest[2]) );
  NOR2X1 U204 ( .A(n83), .B(n182), .Y(neg_dest[3]) );
  NAND3X1 U205 ( .A(n70), .B(instruction_available), .C(n49), .Y(n183) );
  NOR2X1 U206 ( .A(n28), .B(n183), .Y(sin_dest[0]) );
  NOR2X1 U207 ( .A(n68), .B(n183), .Y(sin_dest[1]) );
  NOR2X1 U208 ( .A(n92), .B(n183), .Y(sin_dest[2]) );
  NOR2X1 U209 ( .A(n83), .B(n183), .Y(sin_dest[3]) );
  NAND2X1 U210 ( .A(n67), .B(n218), .Y(n157) );
  NAND2X1 U211 ( .A(N51), .B(n217), .Y(n156) );
  OAI22X1 U212 ( .A(dependency[9]), .B(n157), .C(dependency[10]), .D(n156), 
        .Y(n152) );
  INVX2 U213 ( .A(N52), .Y(n219) );
  NAND2X1 U214 ( .A(n4), .B(n219), .Y(n143) );
  AOI21X1 U215 ( .A(n144), .B(n78), .C(n143), .Y(n145) );
  OAI21X1 U216 ( .A(dependency[8]), .B(n161), .C(n145), .Y(n151) );
  OAI22X1 U217 ( .A(dependency[13]), .B(n53), .C(dependency[14]), .D(n156), 
        .Y(n150) );
  NAND2X1 U218 ( .A(n4), .B(N52), .Y(n146) );
  AOI21X1 U219 ( .A(n78), .B(n147), .C(n146), .Y(n148) );
  OAI21X1 U220 ( .A(dependency[12]), .B(n161), .C(n148), .Y(n149) );
  OAI22X1 U221 ( .A(n152), .B(n151), .C(n150), .D(n149), .Y(n207) );
  OAI22X1 U222 ( .A(n157), .B(dependency[5]), .C(n156), .D(dependency[6]), .Y(
        n165) );
  INVX2 U223 ( .A(N53), .Y(n220) );
  NAND2X1 U224 ( .A(N52), .B(n220), .Y(n153) );
  AOI21X1 U225 ( .A(n78), .B(n154), .C(n153), .Y(n155) );
  OAI21X1 U226 ( .A(dependency[4]), .B(n161), .C(n155), .Y(n164) );
  OAI22X1 U227 ( .A(dependency[1]), .B(n53), .C(n156), .D(dependency[2]), .Y(
        n163) );
  NAND2X1 U228 ( .A(n220), .B(n219), .Y(n158) );
  AOI21X1 U229 ( .A(n78), .B(n159), .C(n158), .Y(n160) );
  OAI21X1 U230 ( .A(n161), .B(dependency[0]), .C(n160), .Y(n162) );
  OAI22X1 U231 ( .A(n165), .B(n164), .C(n163), .D(n162), .Y(n206) );
  NOR2X1 U232 ( .A(n207), .B(n206), .Y(n166) );
  NAND3X1 U233 ( .A(n168), .B(n167), .C(n166), .Y(n169) );
  INVX2 U234 ( .A(n169), .Y(n174) );
  NAND2X1 U235 ( .A(n1), .B(n186), .Y(n172) );
  NOR2X1 U236 ( .A(n172), .B(n171), .Y(n173) );
  NAND3X1 U237 ( .A(n173), .B(n80), .C(n174), .Y(n249) );
  NOR2X1 U238 ( .A(n28), .B(n95), .Y(mul_dest[0]) );
  NOR2X1 U239 ( .A(n68), .B(n95), .Y(mul_dest[1]) );
  NOR2X1 U240 ( .A(n92), .B(n95), .Y(mul_dest[2]) );
  NOR2X1 U241 ( .A(n83), .B(n95), .Y(mul_dest[3]) );
  NAND2X1 U242 ( .A(n1), .B(n6), .Y(n191) );
  NAND2X1 U243 ( .A(n81), .B(n174), .Y(n251) );
  NAND2X1 U244 ( .A(n176), .B(n74), .Y(n184) );
  NOR2X1 U245 ( .A(n28), .B(n184), .Y(sub_dest[0]) );
  NOR2X1 U246 ( .A(n68), .B(n184), .Y(sub_dest[1]) );
  NOR2X1 U247 ( .A(n92), .B(n184), .Y(sub_dest[2]) );
  NOR2X1 U248 ( .A(n83), .B(n184), .Y(sub_dest[3]) );
  NOR2X1 U249 ( .A(instruction1[14]), .B(instruction1[15]), .Y(n177) );
  NAND3X1 U250 ( .A(instruction1[12]), .B(n52), .C(n177), .Y(n192) );
  INVX2 U251 ( .A(n192), .Y(n178) );
  NAND2X1 U252 ( .A(n178), .B(n74), .Y(n223) );
  NOR2X1 U253 ( .A(n28), .B(n223), .Y(add_dest[0]) );
  NOR2X1 U254 ( .A(n68), .B(n223), .Y(add_dest[1]) );
  NOR2X1 U255 ( .A(n92), .B(n223), .Y(add_dest[2]) );
  NOR2X1 U256 ( .A(n83), .B(n223), .Y(add_dest[3]) );
  NOR2X1 U257 ( .A(instruction1[15]), .B(instruction1[12]), .Y(n179) );
  NAND3X1 U258 ( .A(n52), .B(n202), .C(n179), .Y(n193) );
  NAND3X1 U259 ( .A(n180), .B(n80), .C(instruction_available), .Y(n245) );
  NOR2X1 U260 ( .A(n28), .B(n97), .Y(load_dest[0]) );
  NOR2X1 U261 ( .A(n68), .B(n97), .Y(load_dest[1]) );
  NOR2X1 U262 ( .A(n92), .B(n97), .Y(load_dest[2]) );
  NOR2X1 U263 ( .A(n83), .B(n97), .Y(load_dest[3]) );
  INVX2 U264 ( .A(n227), .Y(move_enable) );
  INVX2 U265 ( .A(n181), .Y(abs_enable) );
  INVX2 U266 ( .A(n182), .Y(neg_enable) );
  INVX2 U267 ( .A(n183), .Y(sin_enable) );
  INVX2 U268 ( .A(n184), .Y(sub_enable) );
  INVX2 U269 ( .A(n223), .Y(add_enable) );
  NAND3X1 U270 ( .A(n72), .B(n36), .C(n49), .Y(n240) );
  NAND2X1 U271 ( .A(n186), .B(n202), .Y(n187) );
  NOR2X1 U272 ( .A(n5), .B(n187), .Y(n188) );
  NAND3X1 U273 ( .A(n189), .B(n38), .C(n188), .Y(n239) );
  NAND2X1 U274 ( .A(n80), .B(n190), .Y(n246) );
  NAND2X1 U275 ( .A(n192), .B(n191), .Y(n215) );
  NAND2X1 U276 ( .A(instruction1[12]), .B(n202), .Y(n194) );
  OAI21X1 U277 ( .A(n52), .B(n194), .C(n193), .Y(n198) );
  AOI21X1 U278 ( .A(n19), .B(n59), .C(n196), .Y(n199) );
  NAND3X1 U279 ( .A(n201), .B(n200), .C(n199), .Y(n212) );
  NAND2X1 U280 ( .A(instruction1[15]), .B(n202), .Y(n203) );
  OAI21X1 U281 ( .A(n36), .B(n203), .C(instruction_available), .Y(n211) );
  INVX2 U282 ( .A(n211), .Y(n204) );
  NOR2X1 U283 ( .A(n42), .B(n37), .Y(n205) );
  OAI21X1 U284 ( .A(n57), .B(n55), .C(n205), .Y(n208) );
  NAND2X1 U285 ( .A(n208), .B(n81), .Y(n209) );
  OAI22X1 U286 ( .A(n211), .B(n212), .C(n210), .D(n209), .Y(n213) );
  NAND2X1 U287 ( .A(instruction_available), .B(n215), .Y(n250) );
  OAI21X1 U288 ( .A(n41), .B(n250), .C(n95), .Y(n216) );
  INVX2 U289 ( .A(n216), .Y(n221) );
  NOR2X1 U290 ( .A(n221), .B(n263), .Y(source2[0]) );
  NOR2X1 U291 ( .A(n221), .B(n268), .Y(source2[1]) );
  NOR2X1 U292 ( .A(n221), .B(n269), .Y(source2[2]) );
  NOR2X1 U293 ( .A(n221), .B(n20), .Y(source2[3]) );
  NOR2X1 U294 ( .A(sin_enable), .B(sub_enable), .Y(n222) );
  NAND3X1 U295 ( .A(n223), .B(n95), .C(n222), .Y(n234) );
  NOR2X1 U296 ( .A(n225), .B(n224), .Y(n226) );
  AOI22X1 U297 ( .A(n226), .B(n71), .C(n70), .D(instruction1[12]), .Y(n228) );
  INVX2 U298 ( .A(instruction_available), .Y(n243) );
  OAI21X1 U299 ( .A(n228), .B(n243), .C(n227), .Y(n235) );
  AOI22X1 U300 ( .A(n48), .B(n234), .C(n235), .D(n48), .Y(n230) );
  NAND2X1 U301 ( .A(store2_enable), .B(n43), .Y(n229) );
  NAND2X1 U302 ( .A(n230), .B(n229), .Y(source1[0]) );
  AOI22X1 U303 ( .A(n50), .B(n234), .C(n235), .D(n50), .Y(n232) );
  NAND2X1 U304 ( .A(store2_enable), .B(n90), .Y(n231) );
  NAND2X1 U305 ( .A(n232), .B(n231), .Y(source1[1]) );
  AOI22X1 U306 ( .A(n235), .B(n51), .C(n51), .D(n234), .Y(n233) );
  OAI21X1 U307 ( .A(n92), .B(n239), .C(n233), .Y(source1[2]) );
  AOI22X1 U308 ( .A(n235), .B(n44), .C(n44), .D(n234), .Y(n236) );
  OAI21X1 U309 ( .A(n83), .B(n239), .C(n236), .Y(source1[3]) );
  NOR2X1 U310 ( .A(n263), .B(n97), .Y(sram_address_load[0]) );
  NOR2X1 U311 ( .A(n268), .B(n97), .Y(sram_address_load[1]) );
  NOR2X1 U312 ( .A(n269), .B(n97), .Y(sram_address_load[2]) );
  NOR2X1 U313 ( .A(n20), .B(n97), .Y(sram_address_load[3]) );
  NOR2X1 U314 ( .A(n270), .B(n97), .Y(sram_address_load[4]) );
  NOR2X1 U315 ( .A(n40), .B(n97), .Y(sram_address_load[5]) );
  NOR2X1 U316 ( .A(n271), .B(n97), .Y(sram_address_load[6]) );
  NOR2X1 U317 ( .A(n272), .B(n97), .Y(sram_address_load[7]) );
  OAI22X1 U318 ( .A(n270), .B(n240), .C(n263), .D(n239), .Y(
        sram_address_store[0]) );
  OAI22X1 U319 ( .A(n40), .B(n240), .C(n268), .D(n239), .Y(
        sram_address_store[1]) );
  OAI22X1 U320 ( .A(n271), .B(n240), .C(n269), .D(n239), .Y(
        sram_address_store[2]) );
  OAI22X1 U321 ( .A(n272), .B(n240), .C(n20), .D(n239), .Y(
        sram_address_store[3]) );
  OAI22X1 U322 ( .A(n28), .B(n240), .C(n270), .D(n239), .Y(
        sram_address_store[4]) );
  OAI22X1 U323 ( .A(n68), .B(n240), .C(n40), .D(n239), .Y(
        sram_address_store[5]) );
  OAI22X1 U324 ( .A(n92), .B(n240), .C(n271), .D(n239), .Y(
        sram_address_store[6]) );
  OAI22X1 U325 ( .A(n83), .B(n240), .C(n272), .D(n239), .Y(
        sram_address_store[7]) );
  OAI21X1 U326 ( .A(n243), .B(n242), .C(n241), .Y(n244) );
  NAND3X1 U327 ( .A(n244), .B(n80), .C(n79), .Y(n247) );
  NAND3X1 U328 ( .A(n246), .B(n247), .C(n245), .Y(n248) );
  INVX2 U329 ( .A(n248), .Y(n256) );
  OAI21X1 U330 ( .A(n250), .B(n251), .C(n249), .Y(n252) );
  NOR2X1 U331 ( .A(n33), .B(n253), .Y(dependency_add[0]) );
  NOR2X1 U332 ( .A(n66), .B(n32), .Y(dependency_add[1]) );
  NOR2X1 U333 ( .A(n69), .B(n32), .Y(dependency_add[2]) );
  NOR2X1 U334 ( .A(n260), .B(n253), .Y(dependency_add[3]) );
  NOR2X1 U335 ( .A(n33), .B(n254), .Y(dependency_add[4]) );
  NOR2X1 U336 ( .A(n88), .B(n254), .Y(dependency_add[5]) );
  NOR2X1 U337 ( .A(n69), .B(n254), .Y(dependency_add[6]) );
  NOR2X1 U338 ( .A(n260), .B(n254), .Y(dependency_add[7]) );
  NAND2X1 U339 ( .A(n16), .B(n256), .Y(n258) );
  NOR2X1 U340 ( .A(n64), .B(n257), .Y(dependency_add[8]) );
  NOR2X1 U341 ( .A(n66), .B(n257), .Y(dependency_add[9]) );
  NOR2X1 U342 ( .A(n69), .B(n257), .Y(dependency_add[10]) );
  NOR2X1 U343 ( .A(n260), .B(n257), .Y(dependency_add[11]) );
  NOR2X1 U344 ( .A(n33), .B(n259), .Y(dependency_add[12]) );
  NOR2X1 U345 ( .A(n88), .B(n259), .Y(dependency_add[13]) );
  NOR2X1 U346 ( .A(n69), .B(n27), .Y(dependency_add[14]) );
  NOR2X1 U347 ( .A(n260), .B(n27), .Y(dependency_add[15]) );
endmodule


module flex_indexer_NUM_CNT_BITS4_1 ( clk, n_rst, clear, count_enable, 
        rollover_val, count_out, rollover_flag );
  input [3:0] rollover_val;
  output [3:0] count_out;
  input clk, n_rst, clear, count_enable;
  output rollover_flag;
  wire   n29, n1, n2, n4, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28;
  wire   [3:0] nxt_count;
  assign rollover_flag = 1'b0;

  DFFSR \count_out_reg[0]  ( .D(nxt_count[0]), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(n29) );
  DFFSR \count_out_reg[3]  ( .D(nxt_count[3]), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(count_out[3]) );
  DFFSR \count_out_reg[1]  ( .D(nxt_count[1]), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(count_out[1]) );
  DFFSR \count_out_reg[2]  ( .D(nxt_count[2]), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(count_out[2]) );
  BUFX4 U8 ( .A(count_out[1]), .Y(n1) );
  INVX1 U9 ( .A(count_enable), .Y(n14) );
  INVX2 U10 ( .A(n29), .Y(n2) );
  INVX8 U11 ( .A(n2), .Y(count_out[0]) );
  INVX2 U12 ( .A(clear), .Y(n15) );
  XOR2X1 U13 ( .A(rollover_val[2]), .B(count_out[2]), .Y(n9) );
  XOR2X1 U14 ( .A(rollover_val[1]), .B(n1), .Y(n4) );
  NOR2X1 U15 ( .A(n9), .B(n4), .Y(n12) );
  XNOR2X1 U16 ( .A(count_out[0]), .B(rollover_val[0]), .Y(n11) );
  XNOR2X1 U17 ( .A(count_out[3]), .B(rollover_val[3]), .Y(n10) );
  NAND3X1 U18 ( .A(n12), .B(n11), .C(n10), .Y(n13) );
  NAND3X1 U19 ( .A(n15), .B(n13), .C(count_enable), .Y(n28) );
  INVX2 U20 ( .A(n28), .Y(n24) );
  NAND2X1 U21 ( .A(n24), .B(count_out[0]), .Y(n17) );
  NAND2X1 U22 ( .A(n15), .B(n14), .Y(n27) );
  OAI21X1 U23 ( .A(count_out[0]), .B(n28), .C(n27), .Y(n16) );
  INVX2 U24 ( .A(n16), .Y(n18) );
  MUX2X1 U25 ( .B(n17), .A(n18), .S(n1), .Y(nxt_count[1]) );
  NAND3X1 U26 ( .A(n1), .B(count_out[0]), .C(n24), .Y(n20) );
  OAI21X1 U27 ( .A(n1), .B(n28), .C(n18), .Y(n22) );
  INVX2 U28 ( .A(n22), .Y(n19) );
  MUX2X1 U29 ( .B(n20), .A(n19), .S(count_out[2]), .Y(nxt_count[2]) );
  INVX2 U30 ( .A(n20), .Y(n21) );
  NAND2X1 U31 ( .A(count_out[2]), .B(n21), .Y(n26) );
  INVX2 U32 ( .A(count_out[2]), .Y(n23) );
  AOI21X1 U33 ( .A(n24), .B(n23), .C(n22), .Y(n25) );
  MUX2X1 U34 ( .B(n26), .A(n25), .S(count_out[3]), .Y(nxt_count[3]) );
  MUX2X1 U35 ( .B(n28), .A(n27), .S(count_out[0]), .Y(nxt_count[0]) );
endmodule


module flex_indexer_NUM_CNT_BITS4_0 ( clk, n_rst, clear, count_enable, 
        rollover_val, count_out, rollover_flag );
  input [3:0] rollover_val;
  output [3:0] count_out;
  input clk, n_rst, clear, count_enable;
  output rollover_flag;
  wire   n62, n63, n64, n65, n1, n2, n4, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n22, n24, n25, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57;
  wire   [3:0] nxt_count;
  assign rollover_flag = 1'b0;

  DFFSR \count_out_reg[0]  ( .D(nxt_count[0]), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(n65) );
  DFFSR \count_out_reg[3]  ( .D(nxt_count[3]), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(n62) );
  DFFSR \count_out_reg[1]  ( .D(nxt_count[1]), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(n64) );
  DFFSR \count_out_reg[2]  ( .D(nxt_count[2]), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(n63) );
  INVX1 U8 ( .A(count_out[2]), .Y(n12) );
  INVX1 U9 ( .A(n18), .Y(n4) );
  MUX2X1 U10 ( .B(n56), .A(n57), .S(n32), .Y(nxt_count[0]) );
  INVX2 U11 ( .A(n10), .Y(n32) );
  INVX8 U12 ( .A(n22), .Y(count_out[0]) );
  INVX2 U13 ( .A(n12), .Y(n13) );
  INVX2 U14 ( .A(n16), .Y(n17) );
  INVX4 U15 ( .A(n25), .Y(count_out[2]) );
  NAND2X1 U16 ( .A(n53), .B(n10), .Y(n1) );
  NAND2X1 U17 ( .A(n24), .B(n2), .Y(n37) );
  INVX2 U18 ( .A(n1), .Y(n2) );
  BUFX4 U19 ( .A(n64), .Y(count_out[1]) );
  INVX2 U20 ( .A(n18), .Y(n19) );
  INVX1 U21 ( .A(n47), .Y(n9) );
  INVX1 U22 ( .A(count_out[3]), .Y(n47) );
  BUFX2 U23 ( .A(count_out[0]), .Y(n10) );
  INVX1 U24 ( .A(count_enable), .Y(n11) );
  INVX2 U25 ( .A(count_enable), .Y(n54) );
  NAND2X1 U26 ( .A(n53), .B(n20), .Y(n14) );
  NAND2X1 U27 ( .A(n24), .B(n15), .Y(n43) );
  INVX2 U28 ( .A(n14), .Y(n15) );
  INVX1 U29 ( .A(n13), .Y(n16) );
  INVX1 U30 ( .A(count_out[1]), .Y(n18) );
  AND2X2 U31 ( .A(n19), .B(n10), .Y(n20) );
  INVX1 U32 ( .A(n17), .Y(n39) );
  BUFX4 U33 ( .A(n62), .Y(count_out[3]) );
  INVX2 U34 ( .A(n65), .Y(n22) );
  BUFX2 U35 ( .A(count_enable), .Y(n24) );
  INVX2 U36 ( .A(n63), .Y(n25) );
  INVX1 U37 ( .A(n19), .Y(n45) );
  XOR2X1 U38 ( .A(n47), .B(rollover_val[3]), .Y(n31) );
  XOR2X1 U39 ( .A(n32), .B(rollover_val[0]), .Y(n30) );
  XOR2X1 U40 ( .A(rollover_val[2]), .B(n13), .Y(n28) );
  XOR2X1 U41 ( .A(rollover_val[1]), .B(n4), .Y(n27) );
  NOR2X1 U42 ( .A(n28), .B(n27), .Y(n29) );
  NAND3X1 U43 ( .A(n31), .B(n30), .C(n29), .Y(n33) );
  INVX2 U44 ( .A(clear), .Y(n55) );
  NAND2X1 U45 ( .A(n33), .B(n55), .Y(n38) );
  INVX2 U46 ( .A(n38), .Y(n53) );
  NAND3X1 U47 ( .A(n33), .B(n32), .C(n55), .Y(n48) );
  INVX2 U48 ( .A(n48), .Y(n35) );
  NOR2X1 U49 ( .A(clear), .B(n45), .Y(n34) );
  AOI22X1 U50 ( .A(n19), .B(n35), .C(n54), .D(n34), .Y(n36) );
  OAI21X1 U51 ( .A(n19), .B(n37), .C(n36), .Y(nxt_count[1]) );
  OAI21X1 U52 ( .A(n19), .B(n38), .C(n48), .Y(n41) );
  NOR2X1 U53 ( .A(clear), .B(n39), .Y(n40) );
  AOI22X1 U54 ( .A(n17), .B(n41), .C(n54), .D(n40), .Y(n42) );
  OAI21X1 U55 ( .A(n17), .B(n43), .C(n42), .Y(nxt_count[2]) );
  NAND3X1 U56 ( .A(n17), .B(n20), .C(n47), .Y(n44) );
  OAI21X1 U57 ( .A(n17), .B(n47), .C(n44), .Y(n50) );
  NAND3X1 U58 ( .A(n9), .B(n53), .C(n45), .Y(n46) );
  OAI21X1 U59 ( .A(n48), .B(n47), .C(n46), .Y(n49) );
  AOI21X1 U60 ( .A(n53), .B(n50), .C(n49), .Y(n52) );
  NAND3X1 U61 ( .A(n9), .B(n55), .C(n11), .Y(n51) );
  OAI21X1 U62 ( .A(n52), .B(n11), .C(n51), .Y(nxt_count[3]) );
  NAND2X1 U63 ( .A(n24), .B(n53), .Y(n57) );
  NAND2X1 U64 ( .A(n54), .B(n55), .Y(n56) );
endmodule


module flex_fifo_WIDTH16_DEPTH10_BITS_WIDTH4_BITS_DEPTH4 ( clk, n_rst, 
        r_enable, w_enable, w_data, r_data, full, empty );
  input [15:0] w_data;
  output [15:0] r_data;
  input clk, n_rst, r_enable, w_enable;
  output full, empty;
  wire   n629, _2_net_, \data[9][15] , \data[9][14] , \data[9][13] ,
         \data[9][12] , \data[9][11] , \data[9][10] , \data[9][9] ,
         \data[9][8] , \data[9][7] , \data[9][6] , \data[9][5] , \data[9][4] ,
         \data[9][3] , \data[9][2] , \data[9][1] , \data[9][0] , \data[8][15] ,
         \data[8][14] , \data[8][13] , \data[8][12] , \data[8][11] ,
         \data[8][10] , \data[8][9] , \data[8][8] , \data[8][7] , \data[8][6] ,
         \data[8][5] , \data[8][4] , \data[8][3] , \data[8][2] , \data[8][1] ,
         \data[8][0] , \data[7][15] , \data[7][14] , \data[7][13] ,
         \data[7][12] , \data[7][11] , \data[7][10] , \data[7][9] ,
         \data[7][8] , \data[7][7] , \data[7][6] , \data[7][5] , \data[7][4] ,
         \data[7][3] , \data[7][2] , \data[7][1] , \data[7][0] , \data[6][15] ,
         \data[6][14] , \data[6][13] , \data[6][12] , \data[6][11] ,
         \data[6][10] , \data[6][9] , \data[6][8] , \data[6][7] , \data[6][6] ,
         \data[6][5] , \data[6][4] , \data[6][3] , \data[6][2] , \data[6][1] ,
         \data[6][0] , \data[5][15] , \data[5][14] , \data[5][13] ,
         \data[5][12] , \data[5][11] , \data[5][10] , \data[5][9] ,
         \data[5][8] , \data[5][7] , \data[5][6] , \data[5][5] , \data[5][4] ,
         \data[5][3] , \data[5][2] , \data[5][1] , \data[5][0] , \data[4][15] ,
         \data[4][14] , \data[4][13] , \data[4][12] , \data[4][11] ,
         \data[4][10] , \data[4][9] , \data[4][8] , \data[4][7] , \data[4][6] ,
         \data[4][5] , \data[4][4] , \data[4][3] , \data[4][2] , \data[4][1] ,
         \data[4][0] , \data[3][15] , \data[3][14] , \data[3][13] ,
         \data[3][12] , \data[3][11] , \data[3][10] , \data[3][9] ,
         \data[3][8] , \data[3][7] , \data[3][6] , \data[3][5] , \data[3][4] ,
         \data[3][3] , \data[3][2] , \data[3][1] , \data[3][0] , \data[2][15] ,
         \data[2][14] , \data[2][13] , \data[2][12] , \data[2][11] ,
         \data[2][10] , \data[2][9] , \data[2][8] , \data[2][7] , \data[2][6] ,
         \data[2][5] , \data[2][4] , \data[2][3] , \data[2][2] , \data[2][1] ,
         \data[2][0] , \data[1][15] , \data[1][14] , \data[1][13] ,
         \data[1][12] , \data[1][11] , \data[1][10] , \data[1][9] ,
         \data[1][8] , \data[1][7] , \data[1][6] , \data[1][5] , \data[1][4] ,
         \data[1][3] , \data[1][2] , \data[1][1] , \data[1][0] , \data[0][15] ,
         \data[0][14] , \data[0][13] , \data[0][12] , \data[0][11] ,
         \data[0][10] , \data[0][9] , \data[0][8] , \data[0][7] , \data[0][6] ,
         \data[0][5] , \data[0][4] , \data[0][3] , \data[0][2] , \data[0][1] ,
         \data[0][0] , \nxt_data[9][15] , \nxt_data[9][14] , \nxt_data[9][13] ,
         \nxt_data[9][12] , \nxt_data[9][11] , \nxt_data[9][10] ,
         \nxt_data[9][9] , \nxt_data[9][8] , \nxt_data[9][7] ,
         \nxt_data[9][6] , \nxt_data[9][5] , \nxt_data[9][4] ,
         \nxt_data[9][3] , \nxt_data[9][2] , \nxt_data[9][1] ,
         \nxt_data[9][0] , \nxt_data[8][15] , \nxt_data[8][14] ,
         \nxt_data[8][13] , \nxt_data[8][12] , \nxt_data[8][11] ,
         \nxt_data[8][10] , \nxt_data[8][9] , \nxt_data[8][8] ,
         \nxt_data[8][7] , \nxt_data[8][6] , \nxt_data[8][5] ,
         \nxt_data[8][4] , \nxt_data[8][3] , \nxt_data[8][2] ,
         \nxt_data[8][1] , \nxt_data[8][0] , \nxt_data[7][15] ,
         \nxt_data[7][14] , \nxt_data[7][13] , \nxt_data[7][12] ,
         \nxt_data[7][11] , \nxt_data[7][10] , \nxt_data[7][9] ,
         \nxt_data[7][8] , \nxt_data[7][7] , \nxt_data[7][6] ,
         \nxt_data[7][5] , \nxt_data[7][4] , \nxt_data[7][3] ,
         \nxt_data[7][2] , \nxt_data[7][1] , \nxt_data[7][0] ,
         \nxt_data[6][15] , \nxt_data[6][14] , \nxt_data[6][13] ,
         \nxt_data[6][12] , \nxt_data[6][11] , \nxt_data[6][10] ,
         \nxt_data[6][9] , \nxt_data[6][8] , \nxt_data[6][7] ,
         \nxt_data[6][6] , \nxt_data[6][5] , \nxt_data[6][4] ,
         \nxt_data[6][3] , \nxt_data[6][2] , \nxt_data[6][1] ,
         \nxt_data[6][0] , \nxt_data[5][15] , \nxt_data[5][14] ,
         \nxt_data[5][13] , \nxt_data[5][12] , \nxt_data[5][11] ,
         \nxt_data[5][10] , \nxt_data[5][9] , \nxt_data[5][8] ,
         \nxt_data[5][7] , \nxt_data[5][6] , \nxt_data[5][5] ,
         \nxt_data[5][4] , \nxt_data[5][3] , \nxt_data[5][2] ,
         \nxt_data[5][1] , \nxt_data[5][0] , \nxt_data[4][15] ,
         \nxt_data[4][14] , \nxt_data[4][13] , \nxt_data[4][12] ,
         \nxt_data[4][11] , \nxt_data[4][10] , \nxt_data[4][9] ,
         \nxt_data[4][8] , \nxt_data[4][7] , \nxt_data[4][6] ,
         \nxt_data[4][5] , \nxt_data[4][4] , \nxt_data[4][3] ,
         \nxt_data[4][2] , \nxt_data[4][1] , \nxt_data[4][0] ,
         \nxt_data[3][15] , \nxt_data[3][14] , \nxt_data[3][13] ,
         \nxt_data[3][12] , \nxt_data[3][11] , \nxt_data[3][10] ,
         \nxt_data[3][9] , \nxt_data[3][8] , \nxt_data[3][7] ,
         \nxt_data[3][6] , \nxt_data[3][5] , \nxt_data[3][4] ,
         \nxt_data[3][3] , \nxt_data[3][2] , \nxt_data[3][1] ,
         \nxt_data[3][0] , \nxt_data[2][15] , \nxt_data[2][14] ,
         \nxt_data[2][13] , \nxt_data[2][12] , \nxt_data[2][11] ,
         \nxt_data[2][10] , \nxt_data[2][9] , \nxt_data[2][8] ,
         \nxt_data[2][7] , \nxt_data[2][6] , \nxt_data[2][5] ,
         \nxt_data[2][4] , \nxt_data[2][3] , \nxt_data[2][2] ,
         \nxt_data[2][1] , \nxt_data[2][0] , \nxt_data[1][15] ,
         \nxt_data[1][14] , \nxt_data[1][13] , \nxt_data[1][12] ,
         \nxt_data[1][11] , \nxt_data[1][10] , \nxt_data[1][9] ,
         \nxt_data[1][8] , \nxt_data[1][7] , \nxt_data[1][6] ,
         \nxt_data[1][5] , \nxt_data[1][4] , \nxt_data[1][3] ,
         \nxt_data[1][2] , \nxt_data[1][1] , \nxt_data[1][0] ,
         \nxt_data[0][15] , \nxt_data[0][14] , \nxt_data[0][13] ,
         \nxt_data[0][12] , \nxt_data[0][11] , \nxt_data[0][10] ,
         \nxt_data[0][9] , \nxt_data[0][8] , \nxt_data[0][7] ,
         \nxt_data[0][6] , \nxt_data[0][5] , \nxt_data[0][4] ,
         \nxt_data[0][3] , \nxt_data[0][2] , \nxt_data[0][1] ,
         \nxt_data[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n627;
  wire   [3:0] w_pointer;
  wire   [3:0] r_pointer;

  DFFSR \data_reg[9][15]  ( .D(\nxt_data[9][15] ), .CLK(clk), .R(n270), .S(
        1'b1), .Q(\data[9][15] ) );
  DFFSR \data_reg[9][14]  ( .D(\nxt_data[9][14] ), .CLK(clk), .R(n270), .S(
        1'b1), .Q(\data[9][14] ) );
  DFFSR \data_reg[9][13]  ( .D(\nxt_data[9][13] ), .CLK(clk), .R(n270), .S(
        1'b1), .Q(\data[9][13] ) );
  DFFSR \data_reg[9][12]  ( .D(\nxt_data[9][12] ), .CLK(clk), .R(n270), .S(
        1'b1), .Q(\data[9][12] ) );
  DFFSR \data_reg[9][11]  ( .D(\nxt_data[9][11] ), .CLK(clk), .R(n270), .S(
        1'b1), .Q(\data[9][11] ) );
  DFFSR \data_reg[9][10]  ( .D(\nxt_data[9][10] ), .CLK(clk), .R(n270), .S(
        1'b1), .Q(\data[9][10] ) );
  DFFSR \data_reg[9][9]  ( .D(\nxt_data[9][9] ), .CLK(clk), .R(n270), .S(1'b1), 
        .Q(\data[9][9] ) );
  DFFSR \data_reg[9][8]  ( .D(\nxt_data[9][8] ), .CLK(clk), .R(n270), .S(1'b1), 
        .Q(\data[9][8] ) );
  DFFSR \data_reg[9][7]  ( .D(\nxt_data[9][7] ), .CLK(clk), .R(n270), .S(1'b1), 
        .Q(\data[9][7] ) );
  DFFSR \data_reg[9][6]  ( .D(\nxt_data[9][6] ), .CLK(clk), .R(n270), .S(1'b1), 
        .Q(\data[9][6] ) );
  DFFSR \data_reg[9][5]  ( .D(\nxt_data[9][5] ), .CLK(clk), .R(n270), .S(1'b1), 
        .Q(\data[9][5] ) );
  DFFSR \data_reg[9][4]  ( .D(\nxt_data[9][4] ), .CLK(clk), .R(n270), .S(1'b1), 
        .Q(\data[9][4] ) );
  DFFSR \data_reg[9][3]  ( .D(\nxt_data[9][3] ), .CLK(clk), .R(n269), .S(1'b1), 
        .Q(\data[9][3] ) );
  DFFSR \data_reg[9][2]  ( .D(\nxt_data[9][2] ), .CLK(clk), .R(n269), .S(1'b1), 
        .Q(\data[9][2] ) );
  DFFSR \data_reg[9][1]  ( .D(\nxt_data[9][1] ), .CLK(clk), .R(n269), .S(1'b1), 
        .Q(\data[9][1] ) );
  DFFSR \data_reg[9][0]  ( .D(\nxt_data[9][0] ), .CLK(clk), .R(n269), .S(1'b1), 
        .Q(\data[9][0] ) );
  DFFSR \data_reg[8][15]  ( .D(\nxt_data[8][15] ), .CLK(clk), .R(n269), .S(
        1'b1), .Q(\data[8][15] ) );
  DFFSR \data_reg[8][14]  ( .D(\nxt_data[8][14] ), .CLK(clk), .R(n269), .S(
        1'b1), .Q(\data[8][14] ) );
  DFFSR \data_reg[8][13]  ( .D(\nxt_data[8][13] ), .CLK(clk), .R(n269), .S(
        1'b1), .Q(\data[8][13] ) );
  DFFSR \data_reg[8][12]  ( .D(\nxt_data[8][12] ), .CLK(clk), .R(n269), .S(
        1'b1), .Q(\data[8][12] ) );
  DFFSR \data_reg[8][11]  ( .D(\nxt_data[8][11] ), .CLK(clk), .R(n269), .S(
        1'b1), .Q(\data[8][11] ) );
  DFFSR \data_reg[8][10]  ( .D(\nxt_data[8][10] ), .CLK(clk), .R(n269), .S(
        1'b1), .Q(\data[8][10] ) );
  DFFSR \data_reg[8][9]  ( .D(\nxt_data[8][9] ), .CLK(clk), .R(n269), .S(1'b1), 
        .Q(\data[8][9] ) );
  DFFSR \data_reg[8][8]  ( .D(\nxt_data[8][8] ), .CLK(clk), .R(n269), .S(1'b1), 
        .Q(\data[8][8] ) );
  DFFSR \data_reg[8][7]  ( .D(\nxt_data[8][7] ), .CLK(clk), .R(n269), .S(1'b1), 
        .Q(\data[8][7] ) );
  DFFSR \data_reg[8][6]  ( .D(\nxt_data[8][6] ), .CLK(clk), .R(n268), .S(1'b1), 
        .Q(\data[8][6] ) );
  DFFSR \data_reg[8][5]  ( .D(\nxt_data[8][5] ), .CLK(clk), .R(n268), .S(1'b1), 
        .Q(\data[8][5] ) );
  DFFSR \data_reg[8][4]  ( .D(\nxt_data[8][4] ), .CLK(clk), .R(n268), .S(1'b1), 
        .Q(\data[8][4] ) );
  DFFSR \data_reg[8][3]  ( .D(\nxt_data[8][3] ), .CLK(clk), .R(n268), .S(1'b1), 
        .Q(\data[8][3] ) );
  DFFSR \data_reg[8][2]  ( .D(\nxt_data[8][2] ), .CLK(clk), .R(n268), .S(1'b1), 
        .Q(\data[8][2] ) );
  DFFSR \data_reg[8][1]  ( .D(\nxt_data[8][1] ), .CLK(clk), .R(n268), .S(1'b1), 
        .Q(\data[8][1] ) );
  DFFSR \data_reg[8][0]  ( .D(\nxt_data[8][0] ), .CLK(clk), .R(n268), .S(1'b1), 
        .Q(\data[8][0] ) );
  DFFSR \data_reg[7][15]  ( .D(\nxt_data[7][15] ), .CLK(clk), .R(n268), .S(
        1'b1), .Q(\data[7][15] ) );
  DFFSR \data_reg[7][14]  ( .D(\nxt_data[7][14] ), .CLK(clk), .R(n268), .S(
        1'b1), .Q(\data[7][14] ) );
  DFFSR \data_reg[7][13]  ( .D(\nxt_data[7][13] ), .CLK(clk), .R(n268), .S(
        1'b1), .Q(\data[7][13] ) );
  DFFSR \data_reg[7][12]  ( .D(\nxt_data[7][12] ), .CLK(clk), .R(n268), .S(
        1'b1), .Q(\data[7][12] ) );
  DFFSR \data_reg[7][11]  ( .D(\nxt_data[7][11] ), .CLK(clk), .R(n268), .S(
        1'b1), .Q(\data[7][11] ) );
  DFFSR \data_reg[7][10]  ( .D(\nxt_data[7][10] ), .CLK(clk), .R(n268), .S(
        1'b1), .Q(\data[7][10] ) );
  DFFSR \data_reg[7][9]  ( .D(\nxt_data[7][9] ), .CLK(clk), .R(n267), .S(1'b1), 
        .Q(\data[7][9] ) );
  DFFSR \data_reg[7][8]  ( .D(\nxt_data[7][8] ), .CLK(clk), .R(n267), .S(1'b1), 
        .Q(\data[7][8] ) );
  DFFSR \data_reg[7][7]  ( .D(\nxt_data[7][7] ), .CLK(clk), .R(n267), .S(1'b1), 
        .Q(\data[7][7] ) );
  DFFSR \data_reg[7][6]  ( .D(\nxt_data[7][6] ), .CLK(clk), .R(n267), .S(1'b1), 
        .Q(\data[7][6] ) );
  DFFSR \data_reg[7][5]  ( .D(\nxt_data[7][5] ), .CLK(clk), .R(n267), .S(1'b1), 
        .Q(\data[7][5] ) );
  DFFSR \data_reg[7][4]  ( .D(\nxt_data[7][4] ), .CLK(clk), .R(n267), .S(1'b1), 
        .Q(\data[7][4] ) );
  DFFSR \data_reg[7][3]  ( .D(\nxt_data[7][3] ), .CLK(clk), .R(n267), .S(1'b1), 
        .Q(\data[7][3] ) );
  DFFSR \data_reg[7][2]  ( .D(\nxt_data[7][2] ), .CLK(clk), .R(n267), .S(1'b1), 
        .Q(\data[7][2] ) );
  DFFSR \data_reg[7][1]  ( .D(\nxt_data[7][1] ), .CLK(clk), .R(n267), .S(1'b1), 
        .Q(\data[7][1] ) );
  DFFSR \data_reg[7][0]  ( .D(\nxt_data[7][0] ), .CLK(clk), .R(n267), .S(1'b1), 
        .Q(\data[7][0] ) );
  DFFSR \data_reg[6][15]  ( .D(\nxt_data[6][15] ), .CLK(clk), .R(n267), .S(
        1'b1), .Q(\data[6][15] ) );
  DFFSR \data_reg[6][14]  ( .D(\nxt_data[6][14] ), .CLK(clk), .R(n267), .S(
        1'b1), .Q(\data[6][14] ) );
  DFFSR \data_reg[6][13]  ( .D(\nxt_data[6][13] ), .CLK(clk), .R(n267), .S(
        1'b1), .Q(\data[6][13] ) );
  DFFSR \data_reg[6][12]  ( .D(\nxt_data[6][12] ), .CLK(clk), .R(n266), .S(
        1'b1), .Q(\data[6][12] ) );
  DFFSR \data_reg[6][11]  ( .D(\nxt_data[6][11] ), .CLK(clk), .R(n266), .S(
        1'b1), .Q(\data[6][11] ) );
  DFFSR \data_reg[6][10]  ( .D(\nxt_data[6][10] ), .CLK(clk), .R(n266), .S(
        1'b1), .Q(\data[6][10] ) );
  DFFSR \data_reg[6][9]  ( .D(\nxt_data[6][9] ), .CLK(clk), .R(n266), .S(1'b1), 
        .Q(\data[6][9] ) );
  DFFSR \data_reg[6][8]  ( .D(\nxt_data[6][8] ), .CLK(clk), .R(n266), .S(1'b1), 
        .Q(\data[6][8] ) );
  DFFSR \data_reg[6][7]  ( .D(\nxt_data[6][7] ), .CLK(clk), .R(n266), .S(1'b1), 
        .Q(\data[6][7] ) );
  DFFSR \data_reg[6][6]  ( .D(\nxt_data[6][6] ), .CLK(clk), .R(n266), .S(1'b1), 
        .Q(\data[6][6] ) );
  DFFSR \data_reg[6][5]  ( .D(\nxt_data[6][5] ), .CLK(clk), .R(n266), .S(1'b1), 
        .Q(\data[6][5] ) );
  DFFSR \data_reg[6][4]  ( .D(\nxt_data[6][4] ), .CLK(clk), .R(n266), .S(1'b1), 
        .Q(\data[6][4] ) );
  DFFSR \data_reg[6][3]  ( .D(\nxt_data[6][3] ), .CLK(clk), .R(n266), .S(1'b1), 
        .Q(\data[6][3] ) );
  DFFSR \data_reg[6][2]  ( .D(\nxt_data[6][2] ), .CLK(clk), .R(n266), .S(1'b1), 
        .Q(\data[6][2] ) );
  DFFSR \data_reg[6][1]  ( .D(\nxt_data[6][1] ), .CLK(clk), .R(n266), .S(1'b1), 
        .Q(\data[6][1] ) );
  DFFSR \data_reg[6][0]  ( .D(\nxt_data[6][0] ), .CLK(clk), .R(n266), .S(1'b1), 
        .Q(\data[6][0] ) );
  DFFSR \data_reg[5][15]  ( .D(\nxt_data[5][15] ), .CLK(clk), .R(n265), .S(
        1'b1), .Q(\data[5][15] ) );
  DFFSR \data_reg[5][14]  ( .D(\nxt_data[5][14] ), .CLK(clk), .R(n265), .S(
        1'b1), .Q(\data[5][14] ) );
  DFFSR \data_reg[5][13]  ( .D(\nxt_data[5][13] ), .CLK(clk), .R(n265), .S(
        1'b1), .Q(\data[5][13] ) );
  DFFSR \data_reg[5][12]  ( .D(\nxt_data[5][12] ), .CLK(clk), .R(n265), .S(
        1'b1), .Q(\data[5][12] ) );
  DFFSR \data_reg[5][11]  ( .D(\nxt_data[5][11] ), .CLK(clk), .R(n265), .S(
        1'b1), .Q(\data[5][11] ) );
  DFFSR \data_reg[5][10]  ( .D(\nxt_data[5][10] ), .CLK(clk), .R(n265), .S(
        1'b1), .Q(\data[5][10] ) );
  DFFSR \data_reg[5][9]  ( .D(\nxt_data[5][9] ), .CLK(clk), .R(n265), .S(1'b1), 
        .Q(\data[5][9] ) );
  DFFSR \data_reg[5][8]  ( .D(\nxt_data[5][8] ), .CLK(clk), .R(n265), .S(1'b1), 
        .Q(\data[5][8] ) );
  DFFSR \data_reg[5][7]  ( .D(\nxt_data[5][7] ), .CLK(clk), .R(n265), .S(1'b1), 
        .Q(\data[5][7] ) );
  DFFSR \data_reg[5][6]  ( .D(\nxt_data[5][6] ), .CLK(clk), .R(n265), .S(1'b1), 
        .Q(\data[5][6] ) );
  DFFSR \data_reg[5][5]  ( .D(\nxt_data[5][5] ), .CLK(clk), .R(n265), .S(1'b1), 
        .Q(\data[5][5] ) );
  DFFSR \data_reg[5][4]  ( .D(\nxt_data[5][4] ), .CLK(clk), .R(n265), .S(1'b1), 
        .Q(\data[5][4] ) );
  DFFSR \data_reg[5][3]  ( .D(\nxt_data[5][3] ), .CLK(clk), .R(n265), .S(1'b1), 
        .Q(\data[5][3] ) );
  DFFSR \data_reg[5][2]  ( .D(\nxt_data[5][2] ), .CLK(clk), .R(n264), .S(1'b1), 
        .Q(\data[5][2] ) );
  DFFSR \data_reg[5][1]  ( .D(\nxt_data[5][1] ), .CLK(clk), .R(n264), .S(1'b1), 
        .Q(\data[5][1] ) );
  DFFSR \data_reg[5][0]  ( .D(\nxt_data[5][0] ), .CLK(clk), .R(n264), .S(1'b1), 
        .Q(\data[5][0] ) );
  DFFSR \data_reg[4][15]  ( .D(\nxt_data[4][15] ), .CLK(clk), .R(n264), .S(
        1'b1), .Q(\data[4][15] ) );
  DFFSR \data_reg[4][14]  ( .D(\nxt_data[4][14] ), .CLK(clk), .R(n264), .S(
        1'b1), .Q(\data[4][14] ) );
  DFFSR \data_reg[4][13]  ( .D(\nxt_data[4][13] ), .CLK(clk), .R(n264), .S(
        1'b1), .Q(\data[4][13] ) );
  DFFSR \data_reg[4][12]  ( .D(\nxt_data[4][12] ), .CLK(clk), .R(n264), .S(
        1'b1), .Q(\data[4][12] ) );
  DFFSR \data_reg[4][11]  ( .D(\nxt_data[4][11] ), .CLK(clk), .R(n264), .S(
        1'b1), .Q(\data[4][11] ) );
  DFFSR \data_reg[4][10]  ( .D(\nxt_data[4][10] ), .CLK(clk), .R(n264), .S(
        1'b1), .Q(\data[4][10] ) );
  DFFSR \data_reg[4][9]  ( .D(\nxt_data[4][9] ), .CLK(clk), .R(n264), .S(1'b1), 
        .Q(\data[4][9] ) );
  DFFSR \data_reg[4][8]  ( .D(\nxt_data[4][8] ), .CLK(clk), .R(n264), .S(1'b1), 
        .Q(\data[4][8] ) );
  DFFSR \data_reg[4][7]  ( .D(\nxt_data[4][7] ), .CLK(clk), .R(n264), .S(1'b1), 
        .Q(\data[4][7] ) );
  DFFSR \data_reg[4][6]  ( .D(\nxt_data[4][6] ), .CLK(clk), .R(n264), .S(1'b1), 
        .Q(\data[4][6] ) );
  DFFSR \data_reg[4][5]  ( .D(\nxt_data[4][5] ), .CLK(clk), .R(n263), .S(1'b1), 
        .Q(\data[4][5] ) );
  DFFSR \data_reg[4][4]  ( .D(\nxt_data[4][4] ), .CLK(clk), .R(n263), .S(1'b1), 
        .Q(\data[4][4] ) );
  DFFSR \data_reg[4][3]  ( .D(\nxt_data[4][3] ), .CLK(clk), .R(n263), .S(1'b1), 
        .Q(\data[4][3] ) );
  DFFSR \data_reg[4][2]  ( .D(\nxt_data[4][2] ), .CLK(clk), .R(n263), .S(1'b1), 
        .Q(\data[4][2] ) );
  DFFSR \data_reg[4][1]  ( .D(\nxt_data[4][1] ), .CLK(clk), .R(n263), .S(1'b1), 
        .Q(\data[4][1] ) );
  DFFSR \data_reg[4][0]  ( .D(\nxt_data[4][0] ), .CLK(clk), .R(n263), .S(1'b1), 
        .Q(\data[4][0] ) );
  DFFSR \data_reg[3][15]  ( .D(\nxt_data[3][15] ), .CLK(clk), .R(n263), .S(
        1'b1), .Q(\data[3][15] ) );
  DFFSR \data_reg[3][14]  ( .D(\nxt_data[3][14] ), .CLK(clk), .R(n263), .S(
        1'b1), .Q(\data[3][14] ) );
  DFFSR \data_reg[3][13]  ( .D(\nxt_data[3][13] ), .CLK(clk), .R(n263), .S(
        1'b1), .Q(\data[3][13] ) );
  DFFSR \data_reg[3][12]  ( .D(\nxt_data[3][12] ), .CLK(clk), .R(n263), .S(
        1'b1), .Q(\data[3][12] ) );
  DFFSR \data_reg[3][11]  ( .D(\nxt_data[3][11] ), .CLK(clk), .R(n263), .S(
        1'b1), .Q(\data[3][11] ) );
  DFFSR \data_reg[3][10]  ( .D(\nxt_data[3][10] ), .CLK(clk), .R(n263), .S(
        1'b1), .Q(\data[3][10] ) );
  DFFSR \data_reg[3][9]  ( .D(\nxt_data[3][9] ), .CLK(clk), .R(n263), .S(1'b1), 
        .Q(\data[3][9] ) );
  DFFSR \data_reg[3][8]  ( .D(\nxt_data[3][8] ), .CLK(clk), .R(n262), .S(1'b1), 
        .Q(\data[3][8] ) );
  DFFSR \data_reg[3][7]  ( .D(\nxt_data[3][7] ), .CLK(clk), .R(n262), .S(1'b1), 
        .Q(\data[3][7] ) );
  DFFSR \data_reg[3][6]  ( .D(\nxt_data[3][6] ), .CLK(clk), .R(n262), .S(1'b1), 
        .Q(\data[3][6] ) );
  DFFSR \data_reg[3][5]  ( .D(\nxt_data[3][5] ), .CLK(clk), .R(n262), .S(1'b1), 
        .Q(\data[3][5] ) );
  DFFSR \data_reg[3][4]  ( .D(\nxt_data[3][4] ), .CLK(clk), .R(n262), .S(1'b1), 
        .Q(\data[3][4] ) );
  DFFSR \data_reg[3][3]  ( .D(\nxt_data[3][3] ), .CLK(clk), .R(n262), .S(1'b1), 
        .Q(\data[3][3] ) );
  DFFSR \data_reg[3][2]  ( .D(\nxt_data[3][2] ), .CLK(clk), .R(n262), .S(1'b1), 
        .Q(\data[3][2] ) );
  DFFSR \data_reg[3][1]  ( .D(\nxt_data[3][1] ), .CLK(clk), .R(n262), .S(1'b1), 
        .Q(\data[3][1] ) );
  DFFSR \data_reg[3][0]  ( .D(\nxt_data[3][0] ), .CLK(clk), .R(n262), .S(1'b1), 
        .Q(\data[3][0] ) );
  DFFSR \data_reg[2][15]  ( .D(\nxt_data[2][15] ), .CLK(clk), .R(n262), .S(
        1'b1), .Q(\data[2][15] ) );
  DFFSR \data_reg[2][14]  ( .D(\nxt_data[2][14] ), .CLK(clk), .R(n262), .S(
        1'b1), .Q(\data[2][14] ) );
  DFFSR \data_reg[2][13]  ( .D(\nxt_data[2][13] ), .CLK(clk), .R(n262), .S(
        1'b1), .Q(\data[2][13] ) );
  DFFSR \data_reg[2][12]  ( .D(\nxt_data[2][12] ), .CLK(clk), .R(n262), .S(
        1'b1), .Q(\data[2][12] ) );
  DFFSR \data_reg[2][11]  ( .D(\nxt_data[2][11] ), .CLK(clk), .R(n261), .S(
        1'b1), .Q(\data[2][11] ) );
  DFFSR \data_reg[2][10]  ( .D(\nxt_data[2][10] ), .CLK(clk), .R(n261), .S(
        1'b1), .Q(\data[2][10] ) );
  DFFSR \data_reg[2][9]  ( .D(\nxt_data[2][9] ), .CLK(clk), .R(n261), .S(1'b1), 
        .Q(\data[2][9] ) );
  DFFSR \data_reg[2][8]  ( .D(\nxt_data[2][8] ), .CLK(clk), .R(n261), .S(1'b1), 
        .Q(\data[2][8] ) );
  DFFSR \data_reg[2][7]  ( .D(\nxt_data[2][7] ), .CLK(clk), .R(n261), .S(1'b1), 
        .Q(\data[2][7] ) );
  DFFSR \data_reg[2][6]  ( .D(\nxt_data[2][6] ), .CLK(clk), .R(n261), .S(1'b1), 
        .Q(\data[2][6] ) );
  DFFSR \data_reg[2][5]  ( .D(\nxt_data[2][5] ), .CLK(clk), .R(n261), .S(1'b1), 
        .Q(\data[2][5] ) );
  DFFSR \data_reg[2][4]  ( .D(\nxt_data[2][4] ), .CLK(clk), .R(n261), .S(1'b1), 
        .Q(\data[2][4] ) );
  DFFSR \data_reg[2][3]  ( .D(\nxt_data[2][3] ), .CLK(clk), .R(n261), .S(1'b1), 
        .Q(\data[2][3] ) );
  DFFSR \data_reg[2][2]  ( .D(\nxt_data[2][2] ), .CLK(clk), .R(n261), .S(1'b1), 
        .Q(\data[2][2] ) );
  DFFSR \data_reg[2][1]  ( .D(\nxt_data[2][1] ), .CLK(clk), .R(n261), .S(1'b1), 
        .Q(\data[2][1] ) );
  DFFSR \data_reg[2][0]  ( .D(\nxt_data[2][0] ), .CLK(clk), .R(n261), .S(1'b1), 
        .Q(\data[2][0] ) );
  DFFSR \data_reg[1][15]  ( .D(\nxt_data[1][15] ), .CLK(clk), .R(n261), .S(
        1'b1), .Q(\data[1][15] ) );
  DFFSR \data_reg[1][14]  ( .D(\nxt_data[1][14] ), .CLK(clk), .R(n260), .S(
        1'b1), .Q(\data[1][14] ) );
  DFFSR \data_reg[1][13]  ( .D(\nxt_data[1][13] ), .CLK(clk), .R(n260), .S(
        1'b1), .Q(\data[1][13] ) );
  DFFSR \data_reg[1][12]  ( .D(\nxt_data[1][12] ), .CLK(clk), .R(n260), .S(
        1'b1), .Q(\data[1][12] ) );
  DFFSR \data_reg[1][11]  ( .D(\nxt_data[1][11] ), .CLK(clk), .R(n260), .S(
        1'b1), .Q(\data[1][11] ) );
  DFFSR \data_reg[1][10]  ( .D(\nxt_data[1][10] ), .CLK(clk), .R(n260), .S(
        1'b1), .Q(\data[1][10] ) );
  DFFSR \data_reg[1][9]  ( .D(\nxt_data[1][9] ), .CLK(clk), .R(n260), .S(1'b1), 
        .Q(\data[1][9] ) );
  DFFSR \data_reg[1][8]  ( .D(\nxt_data[1][8] ), .CLK(clk), .R(n260), .S(1'b1), 
        .Q(\data[1][8] ) );
  DFFSR \data_reg[1][7]  ( .D(\nxt_data[1][7] ), .CLK(clk), .R(n260), .S(1'b1), 
        .Q(\data[1][7] ) );
  DFFSR \data_reg[1][6]  ( .D(\nxt_data[1][6] ), .CLK(clk), .R(n260), .S(1'b1), 
        .Q(\data[1][6] ) );
  DFFSR \data_reg[1][5]  ( .D(\nxt_data[1][5] ), .CLK(clk), .R(n260), .S(1'b1), 
        .Q(\data[1][5] ) );
  DFFSR \data_reg[1][4]  ( .D(\nxt_data[1][4] ), .CLK(clk), .R(n260), .S(1'b1), 
        .Q(\data[1][4] ) );
  DFFSR \data_reg[1][3]  ( .D(\nxt_data[1][3] ), .CLK(clk), .R(n260), .S(1'b1), 
        .Q(\data[1][3] ) );
  DFFSR \data_reg[1][2]  ( .D(\nxt_data[1][2] ), .CLK(clk), .R(n260), .S(1'b1), 
        .Q(\data[1][2] ) );
  DFFSR \data_reg[1][1]  ( .D(\nxt_data[1][1] ), .CLK(clk), .R(n259), .S(1'b1), 
        .Q(\data[1][1] ) );
  DFFSR \data_reg[1][0]  ( .D(\nxt_data[1][0] ), .CLK(clk), .R(n259), .S(1'b1), 
        .Q(\data[1][0] ) );
  DFFSR \data_reg[0][15]  ( .D(\nxt_data[0][15] ), .CLK(clk), .R(n259), .S(
        1'b1), .Q(\data[0][15] ) );
  DFFSR \data_reg[0][14]  ( .D(\nxt_data[0][14] ), .CLK(clk), .R(n259), .S(
        1'b1), .Q(\data[0][14] ) );
  DFFSR \data_reg[0][13]  ( .D(\nxt_data[0][13] ), .CLK(clk), .R(n259), .S(
        1'b1), .Q(\data[0][13] ) );
  DFFSR \data_reg[0][12]  ( .D(\nxt_data[0][12] ), .CLK(clk), .R(n259), .S(
        1'b1), .Q(\data[0][12] ) );
  DFFSR \data_reg[0][11]  ( .D(\nxt_data[0][11] ), .CLK(clk), .R(n259), .S(
        1'b1), .Q(\data[0][11] ) );
  DFFSR \data_reg[0][10]  ( .D(\nxt_data[0][10] ), .CLK(clk), .R(n259), .S(
        1'b1), .Q(\data[0][10] ) );
  DFFSR \data_reg[0][9]  ( .D(\nxt_data[0][9] ), .CLK(clk), .R(n259), .S(1'b1), 
        .Q(\data[0][9] ) );
  DFFSR \data_reg[0][8]  ( .D(\nxt_data[0][8] ), .CLK(clk), .R(n259), .S(1'b1), 
        .Q(\data[0][8] ) );
  DFFSR \data_reg[0][7]  ( .D(\nxt_data[0][7] ), .CLK(clk), .R(n259), .S(1'b1), 
        .Q(\data[0][7] ) );
  DFFSR \data_reg[0][6]  ( .D(\nxt_data[0][6] ), .CLK(clk), .R(n259), .S(1'b1), 
        .Q(\data[0][6] ) );
  DFFSR \data_reg[0][5]  ( .D(\nxt_data[0][5] ), .CLK(clk), .R(n259), .S(1'b1), 
        .Q(\data[0][5] ) );
  DFFSR \data_reg[0][4]  ( .D(\nxt_data[0][4] ), .CLK(clk), .R(n258), .S(1'b1), 
        .Q(\data[0][4] ) );
  DFFSR \data_reg[0][3]  ( .D(\nxt_data[0][3] ), .CLK(clk), .R(n258), .S(1'b1), 
        .Q(\data[0][3] ) );
  DFFSR \data_reg[0][2]  ( .D(\nxt_data[0][2] ), .CLK(clk), .R(n258), .S(1'b1), 
        .Q(\data[0][2] ) );
  DFFSR \data_reg[0][1]  ( .D(\nxt_data[0][1] ), .CLK(clk), .R(n258), .S(1'b1), 
        .Q(\data[0][1] ) );
  DFFSR \data_reg[0][0]  ( .D(\nxt_data[0][0] ), .CLK(clk), .R(n258), .S(1'b1), 
        .Q(\data[0][0] ) );
  flex_indexer_NUM_CNT_BITS4_1 Write_pointer ( .clk(clk), .n_rst(n258), 
        .clear(1'b0), .count_enable(n627), .rollover_val({1'b1, 1'b0, 1'b0, 
        1'b1}), .count_out(w_pointer) );
  flex_indexer_NUM_CNT_BITS4_0 Read_pointer ( .clk(clk), .n_rst(n258), .clear(
        1'b0), .count_enable(_2_net_), .rollover_val({1'b1, 1'b0, 1'b0, 1'b1}), 
        .count_out(r_pointer) );
  AND2X2 U6 ( .A(n484), .B(n5), .Y(n1) );
  BUFX4 U164 ( .A(n251), .Y(n2) );
  INVX2 U165 ( .A(r_pointer[1]), .Y(n5) );
  INVX1 U166 ( .A(r_pointer[1]), .Y(n208) );
  INVX4 U167 ( .A(n172), .Y(n255) );
  INVX1 U168 ( .A(n197), .Y(n3) );
  INVX2 U169 ( .A(n240), .Y(n197) );
  BUFX2 U170 ( .A(n209), .Y(n4) );
  INVX4 U171 ( .A(n7), .Y(n6) );
  INVX2 U172 ( .A(n176), .Y(n7) );
  INVX2 U173 ( .A(n7), .Y(n622) );
  INVX2 U174 ( .A(n176), .Y(n412) );
  INVX1 U175 ( .A(n233), .Y(n8) );
  BUFX2 U176 ( .A(n246), .Y(n9) );
  INVX2 U177 ( .A(r_pointer[3]), .Y(n234) );
  INVX1 U178 ( .A(n233), .Y(n241) );
  NAND2X1 U179 ( .A(n177), .B(n1), .Y(n10) );
  INVX2 U180 ( .A(n242), .Y(n254) );
  INVX1 U181 ( .A(n233), .Y(n171) );
  INVX4 U182 ( .A(n233), .Y(n172) );
  INVX1 U183 ( .A(n179), .Y(n173) );
  NAND2X1 U184 ( .A(n172), .B(n174), .Y(n175) );
  NAND2X1 U185 ( .A(n175), .B(n530), .Y(n532) );
  INVX2 U186 ( .A(n531), .Y(n174) );
  INVX4 U187 ( .A(n252), .Y(n201) );
  NOR2X1 U188 ( .A(n228), .B(n208), .Y(n176) );
  INVX2 U189 ( .A(n282), .Y(n627) );
  INVX2 U190 ( .A(n495), .Y(n413) );
  AND2X2 U191 ( .A(n202), .B(n316), .Y(n177) );
  INVX2 U192 ( .A(r_pointer[2]), .Y(n484) );
  AND2X1 U193 ( .A(n225), .B(\data[3][8] ), .Y(n178) );
  INVX1 U194 ( .A(\data[8][10] ), .Y(n513) );
  BUFX2 U195 ( .A(n301), .Y(n179) );
  INVX2 U196 ( .A(n192), .Y(n180) );
  INVX2 U197 ( .A(n285), .Y(n310) );
  INVX1 U198 ( .A(n284), .Y(full) );
  BUFX4 U199 ( .A(n593), .Y(n181) );
  BUFX4 U200 ( .A(n593), .Y(n182) );
  BUFX4 U201 ( .A(n593), .Y(n183) );
  INVX2 U202 ( .A(n305), .Y(n593) );
  BUFX4 U203 ( .A(n592), .Y(n184) );
  BUFX4 U204 ( .A(n592), .Y(n185) );
  BUFX4 U205 ( .A(n592), .Y(n186) );
  INVX2 U206 ( .A(n298), .Y(n592) );
  BUFX4 U207 ( .A(n591), .Y(n187) );
  BUFX4 U208 ( .A(n591), .Y(n188) );
  BUFX4 U209 ( .A(n591), .Y(n189) );
  INVX2 U210 ( .A(n299), .Y(n591) );
  BUFX4 U211 ( .A(n308), .Y(n190) );
  INVX2 U212 ( .A(n190), .Y(n191) );
  BUFX4 U213 ( .A(n311), .Y(n192) );
  BUFX4 U214 ( .A(n597), .Y(n193) );
  BUFX4 U215 ( .A(n597), .Y(n194) );
  BUFX4 U216 ( .A(n597), .Y(n195) );
  INVX2 U217 ( .A(n287), .Y(n597) );
  INVX8 U218 ( .A(n190), .Y(n601) );
  INVX8 U219 ( .A(n192), .Y(n599) );
  INVX2 U220 ( .A(n216), .Y(n217) );
  INVX4 U221 ( .A(n247), .Y(n196) );
  INVX4 U222 ( .A(n247), .Y(n248) );
  INVX2 U223 ( .A(n252), .Y(n203) );
  AND2X2 U224 ( .A(n476), .B(n475), .Y(n215) );
  INVX1 U225 ( .A(n197), .Y(n198) );
  INVX2 U226 ( .A(n248), .Y(n213) );
  INVX2 U227 ( .A(n224), .Y(n199) );
  AND2X1 U228 ( .A(n223), .B(n204), .Y(n226) );
  BUFX4 U229 ( .A(w_pointer[1]), .Y(n200) );
  INVX1 U230 ( .A(n234), .Y(n222) );
  INVX1 U231 ( .A(n319), .Y(n202) );
  NOR2X1 U232 ( .A(r_pointer[1]), .B(r_pointer[2]), .Y(n239) );
  BUFX2 U233 ( .A(n495), .Y(n218) );
  INVX2 U234 ( .A(n5), .Y(n204) );
  INVX1 U235 ( .A(n224), .Y(n227) );
  NAND2X1 U236 ( .A(n172), .B(\data[8][10] ), .Y(n205) );
  NAND2X1 U237 ( .A(n205), .B(n512), .Y(n514) );
  INVX2 U238 ( .A(n629), .Y(n206) );
  INVX4 U239 ( .A(n206), .Y(r_data[15]) );
  INVX2 U240 ( .A(n356), .Y(n209) );
  INVX1 U241 ( .A(n356), .Y(n251) );
  NAND2X1 U242 ( .A(n198), .B(n1), .Y(n210) );
  INVX4 U243 ( .A(n492), .Y(n211) );
  INVX8 U244 ( .A(n211), .Y(n212) );
  NOR2X1 U245 ( .A(r_pointer[3]), .B(r_pointer[0]), .Y(n240) );
  INVX4 U246 ( .A(r_pointer[0]), .Y(n319) );
  BUFX4 U247 ( .A(n204), .Y(n214) );
  NAND2X1 U248 ( .A(n226), .B(n178), .Y(n464) );
  NAND2X1 U249 ( .A(n499), .B(n500), .Y(n216) );
  NAND2X1 U250 ( .A(n217), .B(n498), .Y(r_data[9]) );
  INVX1 U251 ( .A(n251), .Y(n219) );
  INVX4 U252 ( .A(n209), .Y(n252) );
  INVX4 U253 ( .A(n249), .Y(n253) );
  INVX1 U254 ( .A(n212), .Y(n220) );
  INVX4 U255 ( .A(n212), .Y(n608) );
  BUFX4 U256 ( .A(n242), .Y(n221) );
  INVX8 U257 ( .A(n232), .Y(n607) );
  BUFX2 U258 ( .A(r_pointer[0]), .Y(n223) );
  INVX2 U259 ( .A(r_pointer[3]), .Y(n316) );
  INVX4 U260 ( .A(r_pointer[1]), .Y(n224) );
  INVX4 U261 ( .A(n490), .Y(n247) );
  INVX2 U262 ( .A(r_pointer[2]), .Y(n225) );
  NAND2X1 U263 ( .A(n319), .B(n484), .Y(n228) );
  BUFX2 U264 ( .A(n223), .Y(n229) );
  NAND2X1 U265 ( .A(n215), .B(n474), .Y(r_data[8]) );
  INVX1 U266 ( .A(n225), .Y(n230) );
  INVX2 U267 ( .A(n410), .Y(n231) );
  INVX4 U268 ( .A(n231), .Y(n232) );
  INVX8 U269 ( .A(n196), .Y(n613) );
  AND2X2 U270 ( .A(n227), .B(n319), .Y(n244) );
  AND2X2 U271 ( .A(r_pointer[0]), .B(r_pointer[1]), .Y(n243) );
  AND2X2 U272 ( .A(r_pointer[3]), .B(r_pointer[0]), .Y(n242) );
  OR2X2 U273 ( .A(r_pointer[0]), .B(n234), .Y(n233) );
  NAND2X1 U274 ( .A(n1), .B(n9), .Y(n235) );
  NAND2X1 U275 ( .A(n250), .B(n177), .Y(n236) );
  AND2X2 U276 ( .A(n246), .B(n239), .Y(n237) );
  NAND2X1 U277 ( .A(n177), .B(n250), .Y(n238) );
  XNOR2X1 U278 ( .A(n307), .B(n229), .Y(n245) );
  AND2X2 U279 ( .A(r_pointer[0]), .B(n316), .Y(n246) );
  INVX2 U280 ( .A(w_data[0]), .Y(n312) );
  INVX2 U281 ( .A(w_data[1]), .Y(n332) );
  INVX2 U282 ( .A(w_data[2]), .Y(n350) );
  INVX2 U283 ( .A(w_data[3]), .Y(n369) );
  INVX2 U284 ( .A(w_data[4]), .Y(n390) );
  INVX2 U285 ( .A(w_data[5]), .Y(n408) );
  INVX2 U286 ( .A(w_data[6]), .Y(n426) );
  INVX2 U287 ( .A(w_data[7]), .Y(n444) );
  INVX2 U288 ( .A(w_data[8]), .Y(n463) );
  INVX2 U289 ( .A(w_data[9]), .Y(n483) );
  INVX2 U290 ( .A(w_data[10]), .Y(n506) );
  INVX2 U291 ( .A(w_data[11]), .Y(n524) );
  INVX2 U292 ( .A(w_data[12]), .Y(n542) );
  INVX2 U293 ( .A(w_data[13]), .Y(n560) );
  INVX2 U294 ( .A(w_data[14]), .Y(n578) );
  INVX2 U295 ( .A(w_data[15]), .Y(n606) );
  AND2X2 U296 ( .A(n3), .B(n250), .Y(n249) );
  AND2X2 U297 ( .A(n484), .B(n5), .Y(n250) );
  INVX4 U298 ( .A(n611), .Y(n256) );
  INVX4 U299 ( .A(n286), .Y(n605) );
  INVX4 U300 ( .A(n290), .Y(n604) );
  INVX4 U301 ( .A(n293), .Y(n603) );
  INVX4 U302 ( .A(n302), .Y(n595) );
  INVX8 U303 ( .A(n256), .Y(n257) );
  BUFX2 U304 ( .A(n_rst), .Y(n258) );
  BUFX2 U305 ( .A(n_rst), .Y(n259) );
  BUFX2 U306 ( .A(n_rst), .Y(n260) );
  BUFX2 U307 ( .A(n_rst), .Y(n261) );
  BUFX2 U308 ( .A(n_rst), .Y(n262) );
  BUFX2 U309 ( .A(n_rst), .Y(n263) );
  BUFX2 U310 ( .A(n_rst), .Y(n264) );
  BUFX2 U311 ( .A(n_rst), .Y(n265) );
  BUFX2 U312 ( .A(n_rst), .Y(n266) );
  BUFX2 U313 ( .A(n_rst), .Y(n267) );
  BUFX2 U314 ( .A(n_rst), .Y(n268) );
  BUFX2 U315 ( .A(n_rst), .Y(n269) );
  BUFX2 U316 ( .A(n_rst), .Y(n270) );
  INVX2 U317 ( .A(w_pointer[3]), .Y(n295) );
  XOR2X1 U318 ( .A(n295), .B(n222), .Y(n278) );
  INVX2 U319 ( .A(w_pointer[2]), .Y(n296) );
  XOR2X1 U320 ( .A(n296), .B(n230), .Y(n273) );
  INVX2 U321 ( .A(w_pointer[0]), .Y(n307) );
  XOR2X1 U322 ( .A(n214), .B(n200), .Y(n271) );
  NOR2X1 U323 ( .A(n245), .B(n271), .Y(n272) );
  NAND3X1 U324 ( .A(n278), .B(n273), .C(n272), .Y(n283) );
  AND2X2 U325 ( .A(r_enable), .B(n283), .Y(_2_net_) );
  NAND2X1 U326 ( .A(w_pointer[0]), .B(n200), .Y(n274) );
  XOR2X1 U327 ( .A(n173), .B(n273), .Y(n276) );
  INVX2 U328 ( .A(n274), .Y(n301) );
  NAND2X1 U329 ( .A(w_pointer[2]), .B(n301), .Y(n277) );
  OAI21X1 U330 ( .A(n295), .B(n277), .C(n245), .Y(n275) );
  NOR2X1 U331 ( .A(n276), .B(n275), .Y(n281) );
  XNOR2X1 U332 ( .A(n277), .B(n278), .Y(n280) );
  INVX2 U333 ( .A(n200), .Y(n309) );
  FAX1 U334 ( .A(n309), .B(w_pointer[0]), .C(n214), .YS(n279) );
  NAND3X1 U335 ( .A(n281), .B(n280), .C(n279), .Y(n284) );
  NAND2X1 U336 ( .A(w_enable), .B(n284), .Y(n282) );
  INVX2 U337 ( .A(n283), .Y(empty) );
  INVX2 U338 ( .A(\data[7][0] ), .Y(n320) );
  NAND3X1 U339 ( .A(n627), .B(w_pointer[2]), .C(n295), .Y(n285) );
  NAND2X1 U340 ( .A(n310), .B(n179), .Y(n286) );
  MUX2X1 U341 ( .B(n320), .A(n312), .S(n605), .Y(\nxt_data[7][0] ) );
  INVX2 U342 ( .A(\data[4][0] ), .Y(n321) );
  NAND3X1 U343 ( .A(n310), .B(n309), .C(n307), .Y(n287) );
  MUX2X1 U344 ( .B(n321), .A(n312), .S(n193), .Y(\nxt_data[4][0] ) );
  INVX2 U345 ( .A(\data[9][0] ), .Y(n291) );
  NOR2X1 U346 ( .A(n200), .B(w_pointer[2]), .Y(n288) );
  NAND3X1 U347 ( .A(n627), .B(w_pointer[3]), .C(n288), .Y(n289) );
  INVX2 U348 ( .A(n289), .Y(n292) );
  NAND2X1 U349 ( .A(n292), .B(w_pointer[0]), .Y(n290) );
  MUX2X1 U350 ( .B(n291), .A(n312), .S(n604), .Y(\nxt_data[9][0] ) );
  INVX2 U351 ( .A(\data[8][0] ), .Y(n294) );
  NAND2X1 U352 ( .A(n292), .B(n307), .Y(n293) );
  MUX2X1 U353 ( .B(n294), .A(n312), .S(n603), .Y(\nxt_data[8][0] ) );
  INVX2 U354 ( .A(\data[1][0] ), .Y(n318) );
  NAND3X1 U355 ( .A(n627), .B(n296), .C(n295), .Y(n297) );
  INVX2 U356 ( .A(n297), .Y(n304) );
  NAND3X1 U357 ( .A(n304), .B(w_pointer[0]), .C(n309), .Y(n298) );
  MUX2X1 U358 ( .B(n318), .A(n312), .S(n184), .Y(\nxt_data[1][0] ) );
  INVX2 U359 ( .A(\data[0][0] ), .Y(n300) );
  NAND3X1 U360 ( .A(n304), .B(n309), .C(n307), .Y(n299) );
  MUX2X1 U361 ( .B(n300), .A(n312), .S(n187), .Y(\nxt_data[0][0] ) );
  INVX2 U362 ( .A(\data[3][0] ), .Y(n303) );
  NAND2X1 U363 ( .A(n304), .B(n179), .Y(n302) );
  MUX2X1 U364 ( .B(n303), .A(n312), .S(n595), .Y(\nxt_data[3][0] ) );
  INVX2 U365 ( .A(\data[2][0] ), .Y(n306) );
  NAND3X1 U366 ( .A(n304), .B(n200), .C(n307), .Y(n305) );
  MUX2X1 U367 ( .B(n306), .A(n312), .S(n181), .Y(\nxt_data[2][0] ) );
  INVX2 U368 ( .A(\data[6][0] ), .Y(n313) );
  NAND3X1 U369 ( .A(n310), .B(n200), .C(n307), .Y(n308) );
  MUX2X1 U370 ( .B(n313), .A(n312), .S(n601), .Y(\nxt_data[6][0] ) );
  INVX2 U371 ( .A(\data[5][0] ), .Y(n314) );
  NAND3X1 U372 ( .A(n310), .B(w_pointer[0]), .C(n309), .Y(n311) );
  MUX2X1 U373 ( .B(n314), .A(n312), .S(n599), .Y(\nxt_data[5][0] ) );
  NAND2X1 U374 ( .A(n225), .B(n243), .Y(n410) );
  AOI22X1 U375 ( .A(\data[0][0] ), .B(n413), .C(\data[3][0] ), .D(n607), .Y(
        n326) );
  NAND3X1 U376 ( .A(r_pointer[0]), .B(r_pointer[2]), .C(n224), .Y(n356) );
  NAND3X1 U377 ( .A(r_pointer[2]), .B(n319), .C(n199), .Y(n490) );
  OAI22X1 U378 ( .A(n219), .B(n314), .C(n248), .D(n313), .Y(n315) );
  AOI21X1 U379 ( .A(\data[2][0] ), .B(n622), .C(n315), .Y(n325) );
  AOI22X1 U380 ( .A(n221), .B(\data[9][0] ), .C(n172), .D(\data[8][0] ), .Y(
        n317) );
  OAI21X1 U381 ( .A(n238), .B(n318), .C(n317), .Y(n323) );
  NAND3X1 U382 ( .A(r_pointer[2]), .B(n319), .C(n208), .Y(n492) );
  NAND3X1 U383 ( .A(r_pointer[1]), .B(r_pointer[0]), .C(r_pointer[2]), .Y(n611) );
  OAI22X1 U384 ( .A(n212), .B(n321), .C(n257), .D(n320), .Y(n322) );
  NOR2X1 U385 ( .A(n322), .B(n323), .Y(n324) );
  NAND3X1 U386 ( .A(n326), .B(n325), .C(n324), .Y(r_data[0]) );
  INVX2 U387 ( .A(\data[7][1] ), .Y(n338) );
  MUX2X1 U388 ( .B(n338), .A(n332), .S(n605), .Y(\nxt_data[7][1] ) );
  INVX2 U389 ( .A(\data[4][1] ), .Y(n339) );
  MUX2X1 U390 ( .B(n339), .A(n332), .S(n193), .Y(\nxt_data[4][1] ) );
  INVX2 U391 ( .A(\data[9][1] ), .Y(n327) );
  MUX2X1 U392 ( .B(n327), .A(n332), .S(n604), .Y(\nxt_data[9][1] ) );
  INVX2 U393 ( .A(\data[8][1] ), .Y(n328) );
  MUX2X1 U394 ( .B(n328), .A(n332), .S(n603), .Y(\nxt_data[8][1] ) );
  INVX2 U395 ( .A(\data[1][1] ), .Y(n337) );
  MUX2X1 U396 ( .B(n337), .A(n332), .S(n184), .Y(\nxt_data[1][1] ) );
  INVX2 U397 ( .A(\data[0][1] ), .Y(n329) );
  MUX2X1 U398 ( .B(n329), .A(n332), .S(n187), .Y(\nxt_data[0][1] ) );
  INVX2 U399 ( .A(\data[3][1] ), .Y(n330) );
  MUX2X1 U400 ( .B(n330), .A(n332), .S(n595), .Y(\nxt_data[3][1] ) );
  INVX2 U401 ( .A(\data[2][1] ), .Y(n331) );
  MUX2X1 U402 ( .B(n331), .A(n332), .S(n181), .Y(\nxt_data[2][1] ) );
  INVX2 U403 ( .A(\data[6][1] ), .Y(n333) );
  MUX2X1 U404 ( .B(n333), .A(n332), .S(n601), .Y(\nxt_data[6][1] ) );
  INVX2 U405 ( .A(\data[5][1] ), .Y(n334) );
  MUX2X1 U406 ( .B(n334), .A(n332), .S(n599), .Y(\nxt_data[5][1] ) );
  AOI22X1 U407 ( .A(\data[0][1] ), .B(n413), .C(\data[3][1] ), .D(n607), .Y(
        n344) );
  OAI22X1 U408 ( .A(n219), .B(n334), .C(n248), .D(n333), .Y(n335) );
  AOI21X1 U409 ( .A(\data[2][1] ), .B(n622), .C(n335), .Y(n343) );
  AOI22X1 U410 ( .A(\data[9][1] ), .B(n221), .C(\data[8][1] ), .D(n8), .Y(n336) );
  OAI21X1 U411 ( .A(n235), .B(n337), .C(n336), .Y(n341) );
  OAI22X1 U412 ( .A(n212), .B(n339), .C(n257), .D(n338), .Y(n340) );
  NOR2X1 U413 ( .A(n340), .B(n341), .Y(n342) );
  NAND3X1 U414 ( .A(n343), .B(n344), .C(n342), .Y(r_data[1]) );
  INVX2 U415 ( .A(\data[0][2] ), .Y(n351) );
  MUX2X1 U416 ( .B(n351), .A(n350), .S(n187), .Y(\nxt_data[0][2] ) );
  INVX2 U417 ( .A(\data[1][2] ), .Y(n352) );
  MUX2X1 U418 ( .B(n352), .A(n350), .S(n184), .Y(\nxt_data[1][2] ) );
  INVX2 U419 ( .A(\data[2][2] ), .Y(n345) );
  MUX2X1 U420 ( .B(n345), .A(n350), .S(n181), .Y(\nxt_data[2][2] ) );
  INVX2 U421 ( .A(\data[3][2] ), .Y(n346) );
  MUX2X1 U422 ( .B(n346), .A(n350), .S(n595), .Y(\nxt_data[3][2] ) );
  INVX2 U423 ( .A(\data[4][2] ), .Y(n347) );
  MUX2X1 U424 ( .B(n347), .A(n350), .S(n193), .Y(\nxt_data[4][2] ) );
  INVX2 U425 ( .A(\data[5][2] ), .Y(n348) );
  MUX2X1 U426 ( .B(n348), .A(n350), .S(n599), .Y(\nxt_data[5][2] ) );
  INVX2 U427 ( .A(\data[6][2] ), .Y(n349) );
  MUX2X1 U428 ( .B(n349), .A(n350), .S(n601), .Y(\nxt_data[6][2] ) );
  INVX2 U429 ( .A(\data[8][2] ), .Y(n358) );
  MUX2X1 U430 ( .B(n358), .A(n350), .S(n603), .Y(\nxt_data[8][2] ) );
  INVX2 U431 ( .A(\data[9][2] ), .Y(n354) );
  MUX2X1 U432 ( .B(n354), .A(n350), .S(n604), .Y(\nxt_data[9][2] ) );
  INVX2 U433 ( .A(\data[7][2] ), .Y(n355) );
  MUX2X1 U434 ( .B(n355), .A(n350), .S(n605), .Y(\nxt_data[7][2] ) );
  OAI22X1 U435 ( .A(n236), .B(n352), .C(n253), .D(n351), .Y(n353) );
  AOI21X1 U436 ( .A(\data[2][2] ), .B(n6), .C(n353), .Y(n363) );
  AOI22X1 U437 ( .A(\data[3][2] ), .B(n607), .C(\data[4][2] ), .D(n608), .Y(
        n362) );
  OAI22X1 U438 ( .A(n257), .B(n355), .C(n254), .D(n354), .Y(n360) );
  AOI22X1 U439 ( .A(\data[5][2] ), .B(n4), .C(\data[6][2] ), .D(n613), .Y(n357) );
  OAI21X1 U440 ( .A(n255), .B(n358), .C(n357), .Y(n359) );
  NOR2X1 U441 ( .A(n360), .B(n359), .Y(n361) );
  NAND3X1 U442 ( .A(n363), .B(n362), .C(n361), .Y(r_data[2]) );
  INVX2 U443 ( .A(\data[0][3] ), .Y(n370) );
  MUX2X1 U444 ( .B(n370), .A(n369), .S(n187), .Y(\nxt_data[0][3] ) );
  INVX2 U445 ( .A(\data[1][3] ), .Y(n371) );
  MUX2X1 U446 ( .B(n371), .A(n369), .S(n184), .Y(\nxt_data[1][3] ) );
  INVX2 U447 ( .A(\data[2][3] ), .Y(n364) );
  MUX2X1 U448 ( .B(n364), .A(n369), .S(n181), .Y(\nxt_data[2][3] ) );
  INVX2 U449 ( .A(\data[3][3] ), .Y(n365) );
  MUX2X1 U450 ( .B(n365), .A(n369), .S(n595), .Y(\nxt_data[3][3] ) );
  INVX2 U451 ( .A(\data[4][3] ), .Y(n366) );
  MUX2X1 U452 ( .B(n366), .A(n369), .S(n193), .Y(\nxt_data[4][3] ) );
  INVX2 U453 ( .A(\data[5][3] ), .Y(n367) );
  MUX2X1 U454 ( .B(n367), .A(n369), .S(n599), .Y(\nxt_data[5][3] ) );
  INVX2 U455 ( .A(\data[6][3] ), .Y(n368) );
  MUX2X1 U456 ( .B(n368), .A(n369), .S(n601), .Y(\nxt_data[6][3] ) );
  INVX2 U457 ( .A(\data[8][3] ), .Y(n376) );
  MUX2X1 U458 ( .B(n376), .A(n369), .S(n603), .Y(\nxt_data[8][3] ) );
  INVX2 U459 ( .A(\data[9][3] ), .Y(n373) );
  MUX2X1 U460 ( .B(n373), .A(n369), .S(n604), .Y(\nxt_data[9][3] ) );
  INVX2 U461 ( .A(\data[7][3] ), .Y(n374) );
  MUX2X1 U462 ( .B(n374), .A(n369), .S(n605), .Y(\nxt_data[7][3] ) );
  OAI22X1 U463 ( .A(n10), .B(n371), .C(n210), .D(n370), .Y(n372) );
  AOI21X1 U464 ( .A(\data[2][3] ), .B(n6), .C(n372), .Y(n381) );
  AOI22X1 U465 ( .A(\data[3][3] ), .B(n607), .C(\data[4][3] ), .D(n220), .Y(
        n380) );
  OAI22X1 U466 ( .A(n257), .B(n374), .C(n254), .D(n373), .Y(n378) );
  AOI22X1 U467 ( .A(n2), .B(\data[5][3] ), .C(\data[6][3] ), .D(n613), .Y(n375) );
  OAI21X1 U468 ( .A(n255), .B(n376), .C(n375), .Y(n377) );
  NOR2X1 U469 ( .A(n378), .B(n377), .Y(n379) );
  NAND3X1 U470 ( .A(n381), .B(n380), .C(n379), .Y(r_data[3]) );
  INVX2 U471 ( .A(\data[6][4] ), .Y(n382) );
  MUX2X1 U472 ( .B(n382), .A(n390), .S(n601), .Y(\nxt_data[6][4] ) );
  INVX2 U473 ( .A(\data[5][4] ), .Y(n383) );
  MUX2X1 U474 ( .B(n383), .A(n390), .S(n599), .Y(\nxt_data[5][4] ) );
  INVX2 U475 ( .A(\data[7][4] ), .Y(n384) );
  MUX2X1 U476 ( .B(n384), .A(n390), .S(n605), .Y(\nxt_data[7][4] ) );
  INVX2 U477 ( .A(\data[4][4] ), .Y(n385) );
  MUX2X1 U478 ( .B(n385), .A(n390), .S(n193), .Y(\nxt_data[4][4] ) );
  INVX2 U479 ( .A(\data[9][4] ), .Y(n386) );
  MUX2X1 U480 ( .B(n386), .A(n390), .S(n604), .Y(\nxt_data[9][4] ) );
  INVX2 U481 ( .A(\data[8][4] ), .Y(n387) );
  MUX2X1 U482 ( .B(n387), .A(n390), .S(n603), .Y(\nxt_data[8][4] ) );
  INVX2 U483 ( .A(\data[1][4] ), .Y(n388) );
  MUX2X1 U484 ( .B(n388), .A(n390), .S(n184), .Y(\nxt_data[1][4] ) );
  INVX2 U485 ( .A(\data[0][4] ), .Y(n389) );
  MUX2X1 U486 ( .B(n389), .A(n390), .S(n187), .Y(\nxt_data[0][4] ) );
  INVX2 U487 ( .A(\data[3][4] ), .Y(n391) );
  MUX2X1 U488 ( .B(n391), .A(n390), .S(n595), .Y(\nxt_data[3][4] ) );
  INVX2 U489 ( .A(\data[2][4] ), .Y(n392) );
  MUX2X1 U490 ( .B(n392), .A(n390), .S(n181), .Y(\nxt_data[2][4] ) );
  AOI22X1 U491 ( .A(\data[6][4] ), .B(n213), .C(\data[5][4] ), .D(n2), .Y(n399) );
  AOI22X1 U492 ( .A(\data[7][4] ), .B(n256), .C(\data[4][4] ), .D(n608), .Y(
        n398) );
  OAI22X1 U493 ( .A(n412), .B(n392), .C(n232), .D(n391), .Y(n396) );
  AOI22X1 U494 ( .A(\data[9][4] ), .B(n221), .C(n8), .D(\data[8][4] ), .Y(n394) );
  NAND2X1 U495 ( .A(n239), .B(n240), .Y(n495) );
  AOI22X1 U496 ( .A(n237), .B(\data[1][4] ), .C(n413), .D(\data[0][4] ), .Y(
        n393) );
  NAND2X1 U497 ( .A(n394), .B(n393), .Y(n395) );
  NOR2X1 U498 ( .A(n396), .B(n395), .Y(n397) );
  NAND3X1 U499 ( .A(n398), .B(n399), .C(n397), .Y(r_data[4]) );
  INVX2 U500 ( .A(\data[6][5] ), .Y(n400) );
  MUX2X1 U501 ( .B(n400), .A(n408), .S(n601), .Y(\nxt_data[6][5] ) );
  INVX2 U502 ( .A(\data[5][5] ), .Y(n401) );
  MUX2X1 U503 ( .B(n401), .A(n408), .S(n599), .Y(\nxt_data[5][5] ) );
  INVX2 U504 ( .A(\data[7][5] ), .Y(n402) );
  MUX2X1 U505 ( .B(n402), .A(n408), .S(n605), .Y(\nxt_data[7][5] ) );
  INVX2 U506 ( .A(\data[4][5] ), .Y(n403) );
  MUX2X1 U507 ( .B(n403), .A(n408), .S(n193), .Y(\nxt_data[4][5] ) );
  INVX2 U508 ( .A(\data[9][5] ), .Y(n404) );
  MUX2X1 U509 ( .B(n404), .A(n408), .S(n604), .Y(\nxt_data[9][5] ) );
  INVX2 U510 ( .A(\data[8][5] ), .Y(n405) );
  MUX2X1 U511 ( .B(n405), .A(n408), .S(n603), .Y(\nxt_data[8][5] ) );
  INVX2 U512 ( .A(\data[1][5] ), .Y(n406) );
  MUX2X1 U513 ( .B(n406), .A(n408), .S(n184), .Y(\nxt_data[1][5] ) );
  INVX2 U514 ( .A(\data[0][5] ), .Y(n407) );
  MUX2X1 U515 ( .B(n407), .A(n408), .S(n187), .Y(\nxt_data[0][5] ) );
  INVX2 U516 ( .A(\data[3][5] ), .Y(n409) );
  MUX2X1 U517 ( .B(n409), .A(n408), .S(n595), .Y(\nxt_data[3][5] ) );
  INVX2 U518 ( .A(\data[2][5] ), .Y(n411) );
  MUX2X1 U519 ( .B(n411), .A(n408), .S(n181), .Y(\nxt_data[2][5] ) );
  AOI22X1 U520 ( .A(\data[6][5] ), .B(n613), .C(\data[5][5] ), .D(n2), .Y(n420) );
  AOI22X1 U521 ( .A(\data[7][5] ), .B(n256), .C(\data[4][5] ), .D(n608), .Y(
        n419) );
  OAI22X1 U522 ( .A(n412), .B(n411), .C(n232), .D(n409), .Y(n417) );
  AOI22X1 U523 ( .A(n221), .B(\data[9][5] ), .C(n172), .D(\data[8][5] ), .Y(
        n415) );
  AOI22X1 U524 ( .A(n237), .B(\data[1][5] ), .C(n413), .D(\data[0][5] ), .Y(
        n414) );
  NAND2X1 U525 ( .A(n415), .B(n414), .Y(n416) );
  NOR2X1 U526 ( .A(n417), .B(n416), .Y(n418) );
  NAND3X1 U527 ( .A(n420), .B(n419), .C(n418), .Y(r_data[5]) );
  INVX2 U528 ( .A(\data[0][6] ), .Y(n427) );
  MUX2X1 U529 ( .B(n427), .A(n426), .S(n189), .Y(\nxt_data[0][6] ) );
  INVX2 U530 ( .A(\data[1][6] ), .Y(n428) );
  MUX2X1 U531 ( .B(n428), .A(n426), .S(n186), .Y(\nxt_data[1][6] ) );
  INVX2 U532 ( .A(\data[2][6] ), .Y(n421) );
  MUX2X1 U533 ( .B(n421), .A(n426), .S(n183), .Y(\nxt_data[2][6] ) );
  INVX2 U534 ( .A(\data[3][6] ), .Y(n422) );
  MUX2X1 U535 ( .B(n422), .A(n426), .S(n595), .Y(\nxt_data[3][6] ) );
  INVX2 U536 ( .A(\data[4][6] ), .Y(n423) );
  MUX2X1 U537 ( .B(n423), .A(n426), .S(n195), .Y(\nxt_data[4][6] ) );
  INVX2 U538 ( .A(\data[5][6] ), .Y(n424) );
  MUX2X1 U539 ( .B(n424), .A(n426), .S(n599), .Y(\nxt_data[5][6] ) );
  INVX2 U540 ( .A(\data[6][6] ), .Y(n425) );
  MUX2X1 U541 ( .B(n425), .A(n426), .S(n601), .Y(\nxt_data[6][6] ) );
  INVX2 U542 ( .A(\data[8][6] ), .Y(n433) );
  MUX2X1 U543 ( .B(n433), .A(n426), .S(n603), .Y(\nxt_data[8][6] ) );
  INVX2 U544 ( .A(\data[9][6] ), .Y(n430) );
  MUX2X1 U545 ( .B(n430), .A(n426), .S(n604), .Y(\nxt_data[9][6] ) );
  INVX2 U546 ( .A(\data[7][6] ), .Y(n431) );
  MUX2X1 U547 ( .B(n431), .A(n426), .S(n605), .Y(\nxt_data[7][6] ) );
  OAI22X1 U548 ( .A(n10), .B(n428), .C(n253), .D(n427), .Y(n429) );
  AOI21X1 U549 ( .A(\data[2][6] ), .B(n6), .C(n429), .Y(n438) );
  AOI22X1 U550 ( .A(\data[3][6] ), .B(n607), .C(\data[4][6] ), .D(n608), .Y(
        n437) );
  OAI22X1 U551 ( .A(n257), .B(n431), .C(n254), .D(n430), .Y(n435) );
  AOI22X1 U552 ( .A(\data[5][6] ), .B(n4), .C(\data[6][6] ), .D(n613), .Y(n432) );
  OAI21X1 U553 ( .A(n255), .B(n433), .C(n432), .Y(n434) );
  NOR2X1 U554 ( .A(n435), .B(n434), .Y(n436) );
  NAND3X1 U555 ( .A(n437), .B(n438), .C(n436), .Y(r_data[6]) );
  INVX2 U556 ( .A(\data[0][7] ), .Y(n445) );
  MUX2X1 U557 ( .B(n445), .A(n444), .S(n188), .Y(\nxt_data[0][7] ) );
  INVX2 U558 ( .A(\data[1][7] ), .Y(n446) );
  MUX2X1 U559 ( .B(n446), .A(n444), .S(n185), .Y(\nxt_data[1][7] ) );
  INVX2 U560 ( .A(\data[2][7] ), .Y(n439) );
  MUX2X1 U561 ( .B(n439), .A(n444), .S(n182), .Y(\nxt_data[2][7] ) );
  INVX2 U562 ( .A(\data[3][7] ), .Y(n440) );
  MUX2X1 U563 ( .B(n440), .A(n444), .S(n595), .Y(\nxt_data[3][7] ) );
  INVX2 U564 ( .A(\data[4][7] ), .Y(n441) );
  MUX2X1 U565 ( .B(n441), .A(n444), .S(n194), .Y(\nxt_data[4][7] ) );
  INVX2 U566 ( .A(\data[5][7] ), .Y(n442) );
  MUX2X1 U567 ( .B(n442), .A(n444), .S(n599), .Y(\nxt_data[5][7] ) );
  INVX2 U568 ( .A(\data[6][7] ), .Y(n443) );
  MUX2X1 U569 ( .B(n443), .A(n444), .S(n601), .Y(\nxt_data[6][7] ) );
  INVX2 U570 ( .A(\data[8][7] ), .Y(n451) );
  MUX2X1 U571 ( .B(n451), .A(n444), .S(n603), .Y(\nxt_data[8][7] ) );
  INVX2 U572 ( .A(\data[9][7] ), .Y(n448) );
  MUX2X1 U573 ( .B(n448), .A(n444), .S(n604), .Y(\nxt_data[9][7] ) );
  INVX2 U574 ( .A(\data[7][7] ), .Y(n449) );
  MUX2X1 U575 ( .B(n449), .A(n444), .S(n605), .Y(\nxt_data[7][7] ) );
  OAI22X1 U576 ( .A(n235), .B(n446), .C(n253), .D(n445), .Y(n447) );
  AOI21X1 U577 ( .A(\data[2][7] ), .B(n6), .C(n447), .Y(n456) );
  AOI22X1 U578 ( .A(\data[3][7] ), .B(n607), .C(\data[4][7] ), .D(n608), .Y(
        n455) );
  OAI22X1 U579 ( .A(n257), .B(n449), .C(n254), .D(n448), .Y(n453) );
  AOI22X1 U580 ( .A(\data[5][7] ), .B(n203), .C(\data[6][7] ), .D(n613), .Y(
        n450) );
  OAI21X1 U581 ( .A(n255), .B(n451), .C(n450), .Y(n452) );
  NOR2X1 U582 ( .A(n453), .B(n452), .Y(n454) );
  NAND3X1 U583 ( .A(n456), .B(n455), .C(n454), .Y(r_data[7]) );
  INVX2 U584 ( .A(\data[7][8] ), .Y(n457) );
  MUX2X1 U585 ( .B(n457), .A(n463), .S(n605), .Y(\nxt_data[7][8] ) );
  INVX2 U586 ( .A(\data[3][8] ), .Y(n458) );
  MUX2X1 U587 ( .B(n458), .A(n463), .S(n595), .Y(\nxt_data[3][8] ) );
  INVX2 U588 ( .A(\data[2][8] ), .Y(n466) );
  MUX2X1 U589 ( .B(n466), .A(n463), .S(n183), .Y(\nxt_data[2][8] ) );
  INVX2 U590 ( .A(\data[5][8] ), .Y(n459) );
  MUX2X1 U591 ( .B(n459), .A(n463), .S(n599), .Y(\nxt_data[5][8] ) );
  INVX2 U592 ( .A(\data[9][8] ), .Y(n460) );
  MUX2X1 U593 ( .B(n460), .A(n463), .S(n604), .Y(\nxt_data[9][8] ) );
  INVX2 U594 ( .A(\data[8][8] ), .Y(n461) );
  MUX2X1 U595 ( .B(n461), .A(n463), .S(n603), .Y(\nxt_data[8][8] ) );
  INVX2 U596 ( .A(\data[1][8] ), .Y(n462) );
  MUX2X1 U597 ( .B(n462), .A(n463), .S(n186), .Y(\nxt_data[1][8] ) );
  INVX2 U598 ( .A(\data[0][8] ), .Y(n471) );
  MUX2X1 U599 ( .B(n471), .A(n463), .S(n189), .Y(\nxt_data[0][8] ) );
  INVX2 U600 ( .A(\data[6][8] ), .Y(n468) );
  MUX2X1 U601 ( .B(n468), .A(n463), .S(n601), .Y(\nxt_data[6][8] ) );
  INVX2 U602 ( .A(\data[4][8] ), .Y(n469) );
  MUX2X1 U603 ( .B(n469), .A(n463), .S(n195), .Y(\nxt_data[4][8] ) );
  NAND2X1 U604 ( .A(n244), .B(n225), .Y(n465) );
  OAI21X1 U605 ( .A(n466), .B(n465), .C(n464), .Y(n467) );
  AOI21X1 U606 ( .A(\data[7][8] ), .B(n256), .C(n467), .Y(n476) );
  AOI22X1 U607 ( .A(n201), .B(\data[5][8] ), .C(\data[9][8] ), .D(n221), .Y(
        n475) );
  OAI22X1 U608 ( .A(n212), .B(n469), .C(n248), .D(n468), .Y(n473) );
  AOI22X1 U609 ( .A(n241), .B(\data[8][8] ), .C(\data[1][8] ), .D(n237), .Y(
        n470) );
  OAI21X1 U610 ( .A(n471), .B(n218), .C(n470), .Y(n472) );
  NOR2X1 U611 ( .A(n473), .B(n472), .Y(n474) );
  INVX2 U612 ( .A(\data[7][9] ), .Y(n477) );
  MUX2X1 U613 ( .B(n477), .A(n483), .S(n605), .Y(\nxt_data[7][9] ) );
  INVX2 U614 ( .A(\data[3][9] ), .Y(n478) );
  MUX2X1 U615 ( .B(n478), .A(n483), .S(n595), .Y(\nxt_data[3][9] ) );
  INVX2 U616 ( .A(\data[2][9] ), .Y(n487) );
  MUX2X1 U617 ( .B(n487), .A(n483), .S(n182), .Y(\nxt_data[2][9] ) );
  INVX2 U618 ( .A(\data[5][9] ), .Y(n479) );
  MUX2X1 U619 ( .B(n479), .A(n483), .S(n599), .Y(\nxt_data[5][9] ) );
  INVX2 U620 ( .A(\data[9][9] ), .Y(n480) );
  MUX2X1 U621 ( .B(n480), .A(n483), .S(n604), .Y(\nxt_data[9][9] ) );
  INVX2 U622 ( .A(\data[8][9] ), .Y(n481) );
  MUX2X1 U623 ( .B(n481), .A(n483), .S(n603), .Y(\nxt_data[8][9] ) );
  INVX2 U624 ( .A(\data[1][9] ), .Y(n482) );
  MUX2X1 U625 ( .B(n482), .A(n483), .S(n185), .Y(\nxt_data[1][9] ) );
  INVX2 U626 ( .A(\data[0][9] ), .Y(n494) );
  MUX2X1 U627 ( .B(n494), .A(n483), .S(n188), .Y(\nxt_data[0][9] ) );
  INVX2 U628 ( .A(\data[6][9] ), .Y(n489) );
  MUX2X1 U629 ( .B(n489), .A(n483), .S(n601), .Y(\nxt_data[6][9] ) );
  INVX2 U630 ( .A(\data[4][9] ), .Y(n491) );
  MUX2X1 U631 ( .B(n491), .A(n483), .S(n194), .Y(\nxt_data[4][9] ) );
  NAND2X1 U632 ( .A(n244), .B(n225), .Y(n486) );
  NAND3X1 U633 ( .A(n243), .B(n225), .C(\data[3][9] ), .Y(n485) );
  OAI21X1 U634 ( .A(n487), .B(n486), .C(n485), .Y(n488) );
  AOI21X1 U635 ( .A(\data[7][9] ), .B(n256), .C(n488), .Y(n500) );
  AOI22X1 U636 ( .A(n201), .B(\data[5][9] ), .C(\data[9][9] ), .D(n221), .Y(
        n499) );
  OAI22X1 U637 ( .A(n212), .B(n491), .C(n489), .D(n248), .Y(n497) );
  AOI22X1 U638 ( .A(n171), .B(\data[8][9] ), .C(\data[1][9] ), .D(n237), .Y(
        n493) );
  OAI21X1 U639 ( .A(n494), .B(n218), .C(n493), .Y(n496) );
  NOR2X1 U640 ( .A(n497), .B(n496), .Y(n498) );
  INVX2 U641 ( .A(\data[0][10] ), .Y(n507) );
  MUX2X1 U642 ( .B(n507), .A(n506), .S(n189), .Y(\nxt_data[0][10] ) );
  INVX2 U643 ( .A(\data[1][10] ), .Y(n508) );
  MUX2X1 U644 ( .B(n508), .A(n506), .S(n186), .Y(\nxt_data[1][10] ) );
  INVX2 U645 ( .A(\data[2][10] ), .Y(n501) );
  MUX2X1 U646 ( .B(n501), .A(n506), .S(n183), .Y(\nxt_data[2][10] ) );
  INVX2 U647 ( .A(\data[3][10] ), .Y(n502) );
  MUX2X1 U648 ( .B(n502), .A(n506), .S(n595), .Y(\nxt_data[3][10] ) );
  INVX2 U649 ( .A(\data[4][10] ), .Y(n503) );
  MUX2X1 U650 ( .B(n503), .A(n506), .S(n195), .Y(\nxt_data[4][10] ) );
  INVX2 U651 ( .A(\data[5][10] ), .Y(n504) );
  MUX2X1 U652 ( .B(n504), .A(n506), .S(n180), .Y(\nxt_data[5][10] ) );
  INVX2 U653 ( .A(\data[6][10] ), .Y(n505) );
  MUX2X1 U654 ( .B(n505), .A(n506), .S(n601), .Y(\nxt_data[6][10] ) );
  MUX2X1 U655 ( .B(n513), .A(n506), .S(n603), .Y(\nxt_data[8][10] ) );
  INVX2 U656 ( .A(\data[9][10] ), .Y(n510) );
  MUX2X1 U657 ( .B(n510), .A(n506), .S(n604), .Y(\nxt_data[9][10] ) );
  INVX2 U658 ( .A(\data[7][10] ), .Y(n511) );
  MUX2X1 U659 ( .B(n511), .A(n506), .S(n605), .Y(\nxt_data[7][10] ) );
  OAI22X1 U660 ( .A(n236), .B(n508), .C(n253), .D(n507), .Y(n509) );
  AOI21X1 U661 ( .A(\data[2][10] ), .B(n6), .C(n509), .Y(n518) );
  AOI22X1 U662 ( .A(\data[3][10] ), .B(n607), .C(\data[4][10] ), .D(n608), .Y(
        n517) );
  OAI22X1 U663 ( .A(n257), .B(n511), .C(n254), .D(n510), .Y(n515) );
  AOI22X1 U664 ( .A(n2), .B(\data[5][10] ), .C(\data[6][10] ), .D(n613), .Y(
        n512) );
  NOR2X1 U665 ( .A(n515), .B(n514), .Y(n516) );
  NAND3X1 U666 ( .A(n517), .B(n518), .C(n516), .Y(r_data[10]) );
  INVX2 U667 ( .A(\data[0][11] ), .Y(n525) );
  MUX2X1 U668 ( .B(n525), .A(n524), .S(n188), .Y(\nxt_data[0][11] ) );
  INVX2 U669 ( .A(\data[1][11] ), .Y(n526) );
  MUX2X1 U670 ( .B(n526), .A(n524), .S(n185), .Y(\nxt_data[1][11] ) );
  INVX2 U671 ( .A(\data[2][11] ), .Y(n519) );
  MUX2X1 U672 ( .B(n519), .A(n524), .S(n182), .Y(\nxt_data[2][11] ) );
  INVX2 U673 ( .A(\data[3][11] ), .Y(n520) );
  MUX2X1 U674 ( .B(n520), .A(n524), .S(n595), .Y(\nxt_data[3][11] ) );
  INVX2 U675 ( .A(\data[4][11] ), .Y(n521) );
  MUX2X1 U676 ( .B(n521), .A(n524), .S(n194), .Y(\nxt_data[4][11] ) );
  INVX2 U677 ( .A(\data[5][11] ), .Y(n522) );
  MUX2X1 U678 ( .B(n522), .A(n524), .S(n180), .Y(\nxt_data[5][11] ) );
  INVX2 U679 ( .A(\data[6][11] ), .Y(n523) );
  MUX2X1 U680 ( .B(n523), .A(n524), .S(n601), .Y(\nxt_data[6][11] ) );
  INVX2 U681 ( .A(\data[8][11] ), .Y(n531) );
  MUX2X1 U682 ( .B(n531), .A(n524), .S(n603), .Y(\nxt_data[8][11] ) );
  INVX2 U683 ( .A(\data[9][11] ), .Y(n528) );
  MUX2X1 U684 ( .B(n528), .A(n524), .S(n604), .Y(\nxt_data[9][11] ) );
  INVX2 U685 ( .A(\data[7][11] ), .Y(n529) );
  MUX2X1 U686 ( .B(n529), .A(n524), .S(n605), .Y(\nxt_data[7][11] ) );
  OAI22X1 U687 ( .A(n238), .B(n526), .C(n253), .D(n525), .Y(n527) );
  AOI21X1 U688 ( .A(\data[2][11] ), .B(n6), .C(n527), .Y(n536) );
  AOI22X1 U689 ( .A(\data[3][11] ), .B(n607), .C(\data[4][11] ), .D(n608), .Y(
        n535) );
  OAI22X1 U690 ( .A(n257), .B(n529), .C(n254), .D(n528), .Y(n533) );
  AOI22X1 U691 ( .A(\data[5][11] ), .B(n203), .C(\data[6][11] ), .D(n613), .Y(
        n530) );
  NOR2X1 U692 ( .A(n533), .B(n532), .Y(n534) );
  NAND3X1 U693 ( .A(n535), .B(n536), .C(n534), .Y(r_data[11]) );
  INVX2 U694 ( .A(\data[0][12] ), .Y(n543) );
  MUX2X1 U695 ( .B(n543), .A(n542), .S(n189), .Y(\nxt_data[0][12] ) );
  INVX2 U696 ( .A(\data[1][12] ), .Y(n544) );
  MUX2X1 U697 ( .B(n544), .A(n542), .S(n186), .Y(\nxt_data[1][12] ) );
  INVX2 U698 ( .A(\data[2][12] ), .Y(n537) );
  MUX2X1 U699 ( .B(n537), .A(n542), .S(n183), .Y(\nxt_data[2][12] ) );
  INVX2 U700 ( .A(\data[3][12] ), .Y(n538) );
  MUX2X1 U701 ( .B(n538), .A(n542), .S(n595), .Y(\nxt_data[3][12] ) );
  INVX2 U702 ( .A(\data[4][12] ), .Y(n539) );
  MUX2X1 U703 ( .B(n539), .A(n542), .S(n195), .Y(\nxt_data[4][12] ) );
  INVX2 U704 ( .A(\data[5][12] ), .Y(n540) );
  MUX2X1 U705 ( .B(n540), .A(n542), .S(n180), .Y(\nxt_data[5][12] ) );
  INVX2 U706 ( .A(\data[6][12] ), .Y(n541) );
  MUX2X1 U707 ( .B(n541), .A(n542), .S(n601), .Y(\nxt_data[6][12] ) );
  INVX2 U708 ( .A(\data[8][12] ), .Y(n549) );
  MUX2X1 U709 ( .B(n549), .A(n542), .S(n603), .Y(\nxt_data[8][12] ) );
  INVX2 U710 ( .A(\data[9][12] ), .Y(n546) );
  MUX2X1 U711 ( .B(n546), .A(n542), .S(n604), .Y(\nxt_data[9][12] ) );
  INVX2 U712 ( .A(\data[7][12] ), .Y(n547) );
  MUX2X1 U713 ( .B(n547), .A(n542), .S(n605), .Y(\nxt_data[7][12] ) );
  OAI22X1 U714 ( .A(n236), .B(n544), .C(n253), .D(n543), .Y(n545) );
  AOI21X1 U715 ( .A(\data[2][12] ), .B(n6), .C(n545), .Y(n554) );
  AOI22X1 U716 ( .A(\data[3][12] ), .B(n607), .C(\data[4][12] ), .D(n220), .Y(
        n553) );
  OAI22X1 U717 ( .A(n257), .B(n547), .C(n254), .D(n546), .Y(n551) );
  AOI22X1 U718 ( .A(\data[5][12] ), .B(n4), .C(\data[6][12] ), .D(n613), .Y(
        n548) );
  OAI21X1 U719 ( .A(n255), .B(n549), .C(n548), .Y(n550) );
  NOR2X1 U720 ( .A(n551), .B(n550), .Y(n552) );
  NAND3X1 U721 ( .A(n554), .B(n553), .C(n552), .Y(r_data[12]) );
  INVX2 U722 ( .A(\data[0][13] ), .Y(n561) );
  MUX2X1 U723 ( .B(n561), .A(n560), .S(n188), .Y(\nxt_data[0][13] ) );
  INVX2 U724 ( .A(\data[1][13] ), .Y(n562) );
  MUX2X1 U725 ( .B(n562), .A(n560), .S(n185), .Y(\nxt_data[1][13] ) );
  INVX2 U726 ( .A(\data[2][13] ), .Y(n555) );
  MUX2X1 U727 ( .B(n555), .A(n560), .S(n182), .Y(\nxt_data[2][13] ) );
  INVX2 U728 ( .A(\data[3][13] ), .Y(n556) );
  MUX2X1 U729 ( .B(n556), .A(n560), .S(n595), .Y(\nxt_data[3][13] ) );
  INVX2 U730 ( .A(\data[4][13] ), .Y(n557) );
  MUX2X1 U731 ( .B(n557), .A(n560), .S(n194), .Y(\nxt_data[4][13] ) );
  INVX2 U732 ( .A(\data[5][13] ), .Y(n558) );
  MUX2X1 U733 ( .B(n558), .A(n560), .S(n599), .Y(\nxt_data[5][13] ) );
  INVX2 U734 ( .A(\data[6][13] ), .Y(n559) );
  MUX2X1 U735 ( .B(n559), .A(n560), .S(n191), .Y(\nxt_data[6][13] ) );
  INVX2 U736 ( .A(\data[8][13] ), .Y(n567) );
  MUX2X1 U737 ( .B(n567), .A(n560), .S(n603), .Y(\nxt_data[8][13] ) );
  INVX2 U738 ( .A(\data[9][13] ), .Y(n564) );
  MUX2X1 U739 ( .B(n564), .A(n560), .S(n604), .Y(\nxt_data[9][13] ) );
  INVX2 U740 ( .A(\data[7][13] ), .Y(n565) );
  MUX2X1 U741 ( .B(n565), .A(n560), .S(n605), .Y(\nxt_data[7][13] ) );
  OAI22X1 U742 ( .A(n235), .B(n562), .C(n210), .D(n561), .Y(n563) );
  AOI21X1 U743 ( .A(\data[2][13] ), .B(n6), .C(n563), .Y(n572) );
  AOI22X1 U744 ( .A(\data[3][13] ), .B(n607), .C(\data[4][13] ), .D(n608), .Y(
        n571) );
  OAI22X1 U745 ( .A(n257), .B(n565), .C(n254), .D(n564), .Y(n569) );
  AOI22X1 U746 ( .A(\data[5][13] ), .B(n203), .C(\data[6][13] ), .D(n213), .Y(
        n566) );
  OAI21X1 U747 ( .A(n255), .B(n567), .C(n566), .Y(n568) );
  NOR2X1 U748 ( .A(n569), .B(n568), .Y(n570) );
  NAND3X1 U749 ( .A(n572), .B(n571), .C(n570), .Y(r_data[13]) );
  INVX2 U750 ( .A(\data[0][14] ), .Y(n579) );
  MUX2X1 U751 ( .B(n579), .A(n578), .S(n189), .Y(\nxt_data[0][14] ) );
  INVX2 U752 ( .A(\data[1][14] ), .Y(n580) );
  MUX2X1 U753 ( .B(n580), .A(n578), .S(n186), .Y(\nxt_data[1][14] ) );
  INVX2 U754 ( .A(\data[2][14] ), .Y(n573) );
  MUX2X1 U755 ( .B(n573), .A(n578), .S(n183), .Y(\nxt_data[2][14] ) );
  INVX2 U756 ( .A(\data[3][14] ), .Y(n574) );
  MUX2X1 U757 ( .B(n574), .A(n578), .S(n595), .Y(\nxt_data[3][14] ) );
  INVX2 U758 ( .A(\data[4][14] ), .Y(n575) );
  MUX2X1 U759 ( .B(n575), .A(n578), .S(n195), .Y(\nxt_data[4][14] ) );
  INVX2 U760 ( .A(\data[5][14] ), .Y(n576) );
  MUX2X1 U761 ( .B(n576), .A(n578), .S(n599), .Y(\nxt_data[5][14] ) );
  INVX2 U762 ( .A(\data[6][14] ), .Y(n577) );
  MUX2X1 U763 ( .B(n577), .A(n578), .S(n191), .Y(\nxt_data[6][14] ) );
  INVX2 U764 ( .A(\data[8][14] ), .Y(n585) );
  MUX2X1 U765 ( .B(n585), .A(n578), .S(n603), .Y(\nxt_data[8][14] ) );
  INVX2 U766 ( .A(\data[9][14] ), .Y(n582) );
  MUX2X1 U767 ( .B(n582), .A(n578), .S(n604), .Y(\nxt_data[9][14] ) );
  INVX2 U768 ( .A(\data[7][14] ), .Y(n583) );
  MUX2X1 U769 ( .B(n583), .A(n578), .S(n605), .Y(\nxt_data[7][14] ) );
  OAI22X1 U770 ( .A(n236), .B(n580), .C(n210), .D(n579), .Y(n581) );
  AOI21X1 U771 ( .A(\data[2][14] ), .B(n6), .C(n581), .Y(n590) );
  AOI22X1 U772 ( .A(\data[3][14] ), .B(n607), .C(\data[4][14] ), .D(n220), .Y(
        n589) );
  OAI22X1 U773 ( .A(n257), .B(n583), .C(n254), .D(n582), .Y(n587) );
  AOI22X1 U774 ( .A(\data[5][14] ), .B(n2), .C(\data[6][14] ), .D(n213), .Y(
        n584) );
  OAI21X1 U775 ( .A(n255), .B(n585), .C(n584), .Y(n586) );
  NOR2X1 U776 ( .A(n587), .B(n586), .Y(n588) );
  NAND3X1 U777 ( .A(n590), .B(n589), .C(n588), .Y(r_data[14]) );
  INVX2 U778 ( .A(\data[0][15] ), .Y(n619) );
  MUX2X1 U779 ( .B(n619), .A(n606), .S(n188), .Y(\nxt_data[0][15] ) );
  INVX2 U780 ( .A(\data[1][15] ), .Y(n620) );
  MUX2X1 U781 ( .B(n620), .A(n606), .S(n185), .Y(\nxt_data[1][15] ) );
  INVX2 U782 ( .A(\data[2][15] ), .Y(n594) );
  MUX2X1 U783 ( .B(n594), .A(n606), .S(n182), .Y(\nxt_data[2][15] ) );
  INVX2 U784 ( .A(\data[3][15] ), .Y(n596) );
  MUX2X1 U785 ( .B(n596), .A(n606), .S(n595), .Y(\nxt_data[3][15] ) );
  INVX2 U786 ( .A(\data[4][15] ), .Y(n598) );
  MUX2X1 U787 ( .B(n598), .A(n606), .S(n194), .Y(\nxt_data[4][15] ) );
  INVX2 U788 ( .A(\data[5][15] ), .Y(n600) );
  MUX2X1 U789 ( .B(n600), .A(n606), .S(n599), .Y(\nxt_data[5][15] ) );
  INVX2 U790 ( .A(\data[6][15] ), .Y(n602) );
  MUX2X1 U791 ( .B(n602), .A(n606), .S(n191), .Y(\nxt_data[6][15] ) );
  INVX2 U792 ( .A(\data[8][15] ), .Y(n612) );
  MUX2X1 U793 ( .B(n612), .A(n606), .S(n603), .Y(\nxt_data[8][15] ) );
  INVX2 U794 ( .A(\data[9][15] ), .Y(n609) );
  MUX2X1 U795 ( .B(n609), .A(n606), .S(n604), .Y(\nxt_data[9][15] ) );
  INVX2 U796 ( .A(\data[7][15] ), .Y(n610) );
  MUX2X1 U797 ( .B(n610), .A(n606), .S(n605), .Y(\nxt_data[7][15] ) );
  AOI22X1 U798 ( .A(n608), .B(\data[4][15] ), .C(\data[3][15] ), .D(n607), .Y(
        n625) );
  OAI22X1 U799 ( .A(n257), .B(n610), .C(n254), .D(n609), .Y(n618) );
  NOR2X1 U800 ( .A(n255), .B(n612), .Y(n617) );
  NAND2X1 U801 ( .A(\data[5][15] ), .B(n203), .Y(n615) );
  NAND2X1 U802 ( .A(\data[6][15] ), .B(n613), .Y(n614) );
  NAND2X1 U803 ( .A(n615), .B(n614), .Y(n616) );
  NOR3X1 U804 ( .A(n618), .B(n617), .C(n616), .Y(n624) );
  OAI22X1 U805 ( .A(n235), .B(n620), .C(n210), .D(n619), .Y(n621) );
  AOI21X1 U806 ( .A(\data[2][15] ), .B(n6), .C(n621), .Y(n623) );
  NAND3X1 U807 ( .A(n625), .B(n623), .C(n624), .Y(n629) );
endmodule


module dependancy_reg ( clk, n_rst, dependency_set, dependency_remove, 
        dependency_exists );
  input [15:0] dependency_set;
  input [15:0] dependency_remove;
  output [15:0] dependency_exists;
  input clk, n_rst;
  wire   n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n65, n66, n67, n68, n69;

  DFFSR \dependency_exists_reg[15]  ( .D(n64), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(dependency_exists[15]) );
  DFFSR \dependency_exists_reg[14]  ( .D(n63), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(dependency_exists[14]) );
  DFFSR \dependency_exists_reg[13]  ( .D(n62), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(dependency_exists[13]) );
  DFFSR \dependency_exists_reg[12]  ( .D(n61), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(dependency_exists[12]) );
  DFFSR \dependency_exists_reg[11]  ( .D(n60), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(dependency_exists[11]) );
  DFFSR \dependency_exists_reg[10]  ( .D(n59), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(dependency_exists[10]) );
  DFFSR \dependency_exists_reg[9]  ( .D(n58), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(dependency_exists[9]) );
  DFFSR \dependency_exists_reg[8]  ( .D(n57), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(dependency_exists[8]) );
  DFFSR \dependency_exists_reg[7]  ( .D(n56), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(dependency_exists[7]) );
  DFFSR \dependency_exists_reg[6]  ( .D(n55), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(dependency_exists[6]) );
  DFFSR \dependency_exists_reg[5]  ( .D(n54), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(dependency_exists[5]) );
  DFFSR \dependency_exists_reg[4]  ( .D(n53), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(dependency_exists[4]) );
  DFFSR \dependency_exists_reg[3]  ( .D(n52), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(dependency_exists[3]) );
  DFFSR \dependency_exists_reg[2]  ( .D(n51), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(dependency_exists[2]) );
  DFFSR \dependency_exists_reg[1]  ( .D(n50), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(dependency_exists[1]) );
  DFFSR \dependency_exists_reg[0]  ( .D(n49), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(dependency_exists[0]) );
  OR2X2 U19 ( .A(dependency_remove[4]), .B(n31), .Y(n17) );
  NAND2X1 U20 ( .A(n17), .B(n30), .Y(n53) );
  INVX1 U21 ( .A(dependency_exists[4]), .Y(n31) );
  OR2X2 U22 ( .A(dependency_remove[11]), .B(n45), .Y(n18) );
  NAND2X1 U23 ( .A(n18), .B(n44), .Y(n60) );
  INVX1 U24 ( .A(dependency_exists[11]), .Y(n45) );
  OR2X2 U25 ( .A(dependency_remove[7]), .B(n37), .Y(n19) );
  NAND2X1 U26 ( .A(n19), .B(n36), .Y(n56) );
  INVX1 U27 ( .A(dependency_exists[7]), .Y(n37) );
  OR2X2 U28 ( .A(dependency_remove[3]), .B(n29), .Y(n20) );
  NAND2X1 U29 ( .A(n28), .B(n20), .Y(n52) );
  INVX1 U30 ( .A(dependency_exists[3]), .Y(n29) );
  INVX1 U31 ( .A(dependency_set[6]), .Y(n34) );
  OR2X2 U32 ( .A(dependency_remove[15]), .B(n69), .Y(n21) );
  NAND2X1 U33 ( .A(n21), .B(n68), .Y(n64) );
  INVX1 U34 ( .A(dependency_exists[15]), .Y(n69) );
  INVX1 U35 ( .A(dependency_set[7]), .Y(n36) );
  INVX1 U36 ( .A(dependency_set[2]), .Y(n26) );
  INVX1 U37 ( .A(dependency_set[4]), .Y(n30) );
  INVX1 U38 ( .A(dependency_set[3]), .Y(n28) );
  INVX1 U39 ( .A(dependency_set[14]), .Y(n66) );
  INVX1 U40 ( .A(dependency_set[0]), .Y(n22) );
  INVX1 U41 ( .A(dependency_set[1]), .Y(n24) );
  INVX1 U42 ( .A(dependency_set[15]), .Y(n68) );
  INVX1 U43 ( .A(dependency_set[11]), .Y(n44) );
  INVX1 U44 ( .A(dependency_set[12]), .Y(n46) );
  INVX1 U45 ( .A(dependency_set[13]), .Y(n48) );
  INVX1 U46 ( .A(dependency_set[8]), .Y(n38) );
  INVX1 U47 ( .A(dependency_set[5]), .Y(n32) );
  INVX1 U48 ( .A(dependency_set[9]), .Y(n40) );
  INVX1 U49 ( .A(dependency_set[10]), .Y(n42) );
  INVX2 U50 ( .A(dependency_exists[0]), .Y(n23) );
  OAI21X1 U51 ( .A(dependency_remove[0]), .B(n23), .C(n22), .Y(n49) );
  INVX2 U52 ( .A(dependency_exists[1]), .Y(n25) );
  OAI21X1 U53 ( .A(dependency_remove[1]), .B(n25), .C(n24), .Y(n50) );
  INVX2 U54 ( .A(dependency_exists[2]), .Y(n27) );
  OAI21X1 U55 ( .A(dependency_remove[2]), .B(n27), .C(n26), .Y(n51) );
  INVX2 U56 ( .A(dependency_exists[5]), .Y(n33) );
  OAI21X1 U57 ( .A(dependency_remove[5]), .B(n33), .C(n32), .Y(n54) );
  INVX2 U58 ( .A(dependency_exists[6]), .Y(n35) );
  OAI21X1 U59 ( .A(dependency_remove[6]), .B(n35), .C(n34), .Y(n55) );
  INVX2 U60 ( .A(dependency_exists[8]), .Y(n39) );
  OAI21X1 U61 ( .A(dependency_remove[8]), .B(n39), .C(n38), .Y(n57) );
  INVX2 U62 ( .A(dependency_exists[9]), .Y(n41) );
  OAI21X1 U63 ( .A(dependency_remove[9]), .B(n41), .C(n40), .Y(n58) );
  INVX2 U64 ( .A(dependency_exists[10]), .Y(n43) );
  OAI21X1 U65 ( .A(dependency_remove[10]), .B(n43), .C(n42), .Y(n59) );
  INVX2 U66 ( .A(dependency_exists[12]), .Y(n47) );
  OAI21X1 U67 ( .A(dependency_remove[12]), .B(n47), .C(n46), .Y(n61) );
  INVX2 U68 ( .A(dependency_exists[13]), .Y(n65) );
  OAI21X1 U69 ( .A(dependency_remove[13]), .B(n65), .C(n48), .Y(n62) );
  INVX2 U70 ( .A(dependency_exists[14]), .Y(n67) );
  OAI21X1 U71 ( .A(dependency_remove[14]), .B(n67), .C(n66), .Y(n63) );
endmodule


module scheduler ( n_rst, clk, instruction, add_instruction, drop_dependency, 
        buffer_full, sram_address_store, sram_address_load, source1, source2, 
        store2_enable, store1_enable, load_enable, add_enable, sub_enable, 
        mul_enable, sin_enable, neg_enable, abs_enable, move_enable, load_dest, 
        add_dest, sub_dest, mul_dest, sin_dest, neg_dest, abs_dest, move_dest
 );
  input [15:0] instruction;
  input [15:0] drop_dependency;
  output [7:0] sram_address_store;
  output [7:0] sram_address_load;
  output [3:0] source1;
  output [3:0] source2;
  output [3:0] load_dest;
  output [3:0] add_dest;
  output [3:0] sub_dest;
  output [3:0] mul_dest;
  output [3:0] sin_dest;
  output [3:0] neg_dest;
  output [3:0] abs_dest;
  output [3:0] move_dest;
  input n_rst, clk, add_instruction;
  output buffer_full, store2_enable, store1_enable, load_enable, add_enable,
         sub_enable, mul_enable, sin_enable, neg_enable, abs_enable,
         move_enable;
  wire   buff_read_enable, empty, n2, n3, n4;
  wire   [15:0] buffer_head;
  wire   [15:0] curr_dependents;
  wire   [15:0] dependnecy_add;

  scheduling_logic Logic ( .instruction1({buffer_head[15:13], n3, 
        buffer_head[11:0]}), .dependency(curr_dependents), 
        .instruction_available(n4), .dependency_add(dependnecy_add), 
        .sram_address_store(sram_address_store), .sram_address_load(
        sram_address_load), .source1(source1), .source2(source2), 
        .read_instruction1(buff_read_enable), .store2_enable(store2_enable), 
        .store1_enable(store1_enable), .load_enable(load_enable), .add_enable(
        add_enable), .sub_enable(sub_enable), .mul_enable(mul_enable), 
        .sin_enable(sin_enable), .neg_enable(neg_enable), .abs_enable(
        abs_enable), .move_enable(move_enable), .load_dest(load_dest), 
        .add_dest(add_dest), .sub_dest(sub_dest), .mul_dest(mul_dest), 
        .sin_dest(sin_dest), .neg_dest(neg_dest), .abs_dest(abs_dest), 
        .move_dest(move_dest) );
  flex_fifo_WIDTH16_DEPTH10_BITS_WIDTH4_BITS_DEPTH4 Input_Buffer ( .clk(clk), 
        .n_rst(n_rst), .r_enable(buff_read_enable), .w_enable(add_instruction), 
        .w_data(instruction), .r_data(buffer_head), .full(buffer_full), 
        .empty(empty) );
  dependancy_reg Dependency_reg ( .clk(clk), .n_rst(n_rst), .dependency_set(
        dependnecy_add), .dependency_remove(drop_dependency), 
        .dependency_exists(curr_dependents) );
  INVX2 U2 ( .A(buffer_head[12]), .Y(n2) );
  INVX4 U3 ( .A(n2), .Y(n3) );
  INVX2 U4 ( .A(empty), .Y(n4) );
endmodule

