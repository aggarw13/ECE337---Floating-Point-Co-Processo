
module dependency_remove ( .result_address({\result_address[5][3] , 
        \result_address[5][2] , \result_address[5][1] , \result_address[5][0] , 
        \result_address[4][3] , \result_address[4][2] , \result_address[4][1] , 
        \result_address[4][0] , \result_address[3][3] , \result_address[3][2] , 
        \result_address[3][1] , \result_address[3][0] , \result_address[2][3] , 
        \result_address[2][2] , \result_address[2][1] , \result_address[2][0] , 
        \result_address[1][3] , \result_address[1][2] , \result_address[1][1] , 
        \result_address[1][0] , \result_address[0][3] , \result_address[0][2] , 
        \result_address[0][1] , \result_address[0][0] }), remove_enable, 
        dependency_remove );
  input [5:0] remove_enable;
  output [15:0] dependency_remove;
  input \result_address[5][3] , \result_address[5][2] , \result_address[5][1] ,
         \result_address[5][0] , \result_address[4][3] ,
         \result_address[4][2] , \result_address[4][1] ,
         \result_address[4][0] , \result_address[3][3] ,
         \result_address[3][2] , \result_address[3][1] ,
         \result_address[3][0] , \result_address[2][3] ,
         \result_address[2][2] , \result_address[2][1] ,
         \result_address[2][0] , \result_address[1][3] ,
         \result_address[1][2] , \result_address[1][1] ,
         \result_address[1][0] , \result_address[0][3] ,
         \result_address[0][2] , \result_address[0][1] ,
         \result_address[0][0] ;
  wire   n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300;

  OR2X1 U167 ( .A(n149), .B(n150), .Y(dependency_remove[9]) );
  OAI21X1 U168 ( .A(n151), .B(n152), .C(n153), .Y(n150) );
  AOI22X1 U169 ( .A(n154), .B(n155), .C(n156), .D(n157), .Y(n153) );
  OAI21X1 U170 ( .A(n158), .B(n159), .C(n160), .Y(n149) );
  AOI22X1 U171 ( .A(n161), .B(n162), .C(n163), .D(n164), .Y(n160) );
  OR2X1 U172 ( .A(n165), .B(n166), .Y(dependency_remove[8]) );
  OAI21X1 U173 ( .A(n152), .B(n167), .C(n168), .Y(n166) );
  AOI22X1 U174 ( .A(n169), .B(n155), .C(n170), .D(n157), .Y(n168) );
  OAI21X1 U175 ( .A(n159), .B(n171), .C(n172), .Y(n165) );
  AOI22X1 U176 ( .A(n173), .B(n162), .C(n174), .D(n164), .Y(n172) );
  OR2X1 U177 ( .A(n175), .B(n176), .Y(dependency_remove[7]) );
  OAI21X1 U178 ( .A(n177), .B(n178), .C(n179), .Y(n176) );
  AOI22X1 U179 ( .A(n180), .B(n181), .C(n182), .D(n183), .Y(n179) );
  OAI21X1 U180 ( .A(n184), .B(n185), .C(n186), .Y(n175) );
  AOI22X1 U181 ( .A(n187), .B(n188), .C(n189), .D(n190), .Y(n186) );
  OR2X1 U182 ( .A(n191), .B(n192), .Y(dependency_remove[6]) );
  OAI21X1 U183 ( .A(n178), .B(n193), .C(n194), .Y(n192) );
  AOI22X1 U184 ( .A(n195), .B(n181), .C(n196), .D(n183), .Y(n194) );
  OAI21X1 U185 ( .A(n185), .B(n197), .C(n198), .Y(n191) );
  AOI22X1 U186 ( .A(n199), .B(n188), .C(n200), .D(n190), .Y(n198) );
  OR2X1 U187 ( .A(n201), .B(n202), .Y(dependency_remove[5]) );
  OAI21X1 U188 ( .A(n177), .B(n203), .C(n204), .Y(n202) );
  AOI22X1 U189 ( .A(n205), .B(n180), .C(n206), .D(n182), .Y(n204) );
  OAI21X1 U190 ( .A(n184), .B(n207), .C(n208), .Y(n201) );
  AOI22X1 U191 ( .A(n209), .B(n187), .C(n210), .D(n189), .Y(n208) );
  OR2X1 U192 ( .A(n211), .B(n212), .Y(dependency_remove[4]) );
  OAI21X1 U193 ( .A(n193), .B(n203), .C(n213), .Y(n212) );
  AOI22X1 U194 ( .A(n205), .B(n195), .C(n206), .D(n196), .Y(n213) );
  OAI21X1 U195 ( .A(n197), .B(n207), .C(n214), .Y(n211) );
  AOI22X1 U196 ( .A(n209), .B(n199), .C(n210), .D(n200), .Y(n214) );
  OR2X1 U197 ( .A(n215), .B(n216), .Y(dependency_remove[3]) );
  OAI21X1 U198 ( .A(n177), .B(n217), .C(n218), .Y(n216) );
  AOI22X1 U199 ( .A(n219), .B(n180), .C(n220), .D(n182), .Y(n218) );
  OAI21X1 U200 ( .A(n184), .B(n221), .C(n222), .Y(n215) );
  AOI22X1 U201 ( .A(n223), .B(n187), .C(n224), .D(n189), .Y(n222) );
  OR2X1 U202 ( .A(n225), .B(n226), .Y(dependency_remove[2]) );
  OAI21X1 U203 ( .A(n193), .B(n217), .C(n227), .Y(n226) );
  AOI22X1 U204 ( .A(n219), .B(n195), .C(n220), .D(n196), .Y(n227) );
  OAI21X1 U205 ( .A(n197), .B(n221), .C(n228), .Y(n225) );
  AOI22X1 U206 ( .A(n223), .B(n199), .C(n224), .D(n200), .Y(n228) );
  OR2X1 U207 ( .A(n229), .B(n230), .Y(dependency_remove[1]) );
  OAI21X1 U208 ( .A(n152), .B(n177), .C(n231), .Y(n230) );
  AOI22X1 U209 ( .A(n180), .B(n155), .C(n182), .D(n157), .Y(n231) );
  INVX1 U210 ( .A(n232), .Y(n182) );
  NAND3X1 U211 ( .A(remove_enable[4]), .B(n233), .C(\result_address[4][0] ), 
        .Y(n232) );
  INVX1 U212 ( .A(n234), .Y(n180) );
  NAND3X1 U213 ( .A(remove_enable[3]), .B(n235), .C(\result_address[3][0] ), 
        .Y(n234) );
  NAND3X1 U214 ( .A(remove_enable[5]), .B(n236), .C(\result_address[5][0] ), 
        .Y(n177) );
  OAI21X1 U215 ( .A(n159), .B(n184), .C(n237), .Y(n229) );
  AOI22X1 U216 ( .A(n187), .B(n162), .C(n189), .D(n164), .Y(n237) );
  INVX1 U217 ( .A(n238), .Y(n189) );
  NAND3X1 U218 ( .A(remove_enable[1]), .B(n239), .C(\result_address[1][0] ), 
        .Y(n238) );
  INVX1 U219 ( .A(n240), .Y(n187) );
  NAND3X1 U220 ( .A(remove_enable[0]), .B(n241), .C(\result_address[0][0] ), 
        .Y(n240) );
  NAND3X1 U221 ( .A(remove_enable[2]), .B(n242), .C(\result_address[2][0] ), 
        .Y(n184) );
  OR2X1 U222 ( .A(n243), .B(n244), .Y(dependency_remove[15]) );
  OAI21X1 U223 ( .A(n151), .B(n178), .C(n245), .Y(n244) );
  AOI22X1 U224 ( .A(n181), .B(n154), .C(n183), .D(n156), .Y(n245) );
  OAI21X1 U225 ( .A(n158), .B(n185), .C(n246), .Y(n243) );
  AOI22X1 U226 ( .A(n188), .B(n161), .C(n190), .D(n163), .Y(n246) );
  OR2X1 U227 ( .A(n247), .B(n248), .Y(dependency_remove[14]) );
  OAI21X1 U228 ( .A(n167), .B(n178), .C(n249), .Y(n248) );
  AOI22X1 U229 ( .A(n181), .B(n169), .C(n183), .D(n170), .Y(n249) );
  NOR2X1 U230 ( .A(n250), .B(n251), .Y(n183) );
  NOR2X1 U231 ( .A(n252), .B(n253), .Y(n181) );
  NAND2X1 U232 ( .A(\result_address[5][2] ), .B(\result_address[5][1] ), .Y(
        n178) );
  OAI21X1 U233 ( .A(n171), .B(n185), .C(n254), .Y(n247) );
  AOI22X1 U234 ( .A(n188), .B(n173), .C(n190), .D(n174), .Y(n254) );
  NOR2X1 U235 ( .A(n255), .B(n256), .Y(n190) );
  NOR2X1 U236 ( .A(n257), .B(n258), .Y(n188) );
  NAND2X1 U237 ( .A(\result_address[2][2] ), .B(\result_address[2][1] ), .Y(
        n185) );
  OR2X1 U238 ( .A(n259), .B(n260), .Y(dependency_remove[13]) );
  OAI21X1 U239 ( .A(n151), .B(n203), .C(n261), .Y(n260) );
  AOI22X1 U240 ( .A(n205), .B(n154), .C(n206), .D(n156), .Y(n261) );
  OAI21X1 U241 ( .A(n158), .B(n207), .C(n262), .Y(n259) );
  AOI22X1 U242 ( .A(n209), .B(n161), .C(n210), .D(n163), .Y(n262) );
  OR2X1 U243 ( .A(n263), .B(n264), .Y(dependency_remove[12]) );
  OAI21X1 U244 ( .A(n167), .B(n203), .C(n265), .Y(n264) );
  AOI22X1 U245 ( .A(n205), .B(n169), .C(n206), .D(n170), .Y(n265) );
  NOR2X1 U246 ( .A(n250), .B(\result_address[4][1] ), .Y(n206) );
  INVX1 U247 ( .A(\result_address[4][2] ), .Y(n250) );
  NOR2X1 U248 ( .A(n252), .B(\result_address[3][1] ), .Y(n205) );
  INVX1 U249 ( .A(\result_address[3][2] ), .Y(n252) );
  NAND2X1 U250 ( .A(\result_address[5][2] ), .B(n266), .Y(n203) );
  OAI21X1 U251 ( .A(n171), .B(n207), .C(n267), .Y(n263) );
  AOI22X1 U252 ( .A(n209), .B(n173), .C(n210), .D(n174), .Y(n267) );
  NOR2X1 U253 ( .A(n255), .B(\result_address[1][1] ), .Y(n210) );
  INVX1 U254 ( .A(\result_address[1][2] ), .Y(n255) );
  NOR2X1 U255 ( .A(n257), .B(\result_address[0][1] ), .Y(n209) );
  INVX1 U256 ( .A(\result_address[0][2] ), .Y(n257) );
  NAND2X1 U257 ( .A(\result_address[2][2] ), .B(n268), .Y(n207) );
  OR2X1 U258 ( .A(n269), .B(n270), .Y(dependency_remove[11]) );
  OAI21X1 U259 ( .A(n151), .B(n217), .C(n271), .Y(n270) );
  AOI22X1 U260 ( .A(n219), .B(n154), .C(n220), .D(n156), .Y(n271) );
  INVX1 U261 ( .A(n272), .Y(n156) );
  NAND3X1 U262 ( .A(\result_address[4][0] ), .B(remove_enable[4]), .C(
        \result_address[4][3] ), .Y(n272) );
  INVX1 U263 ( .A(n273), .Y(n154) );
  NAND3X1 U264 ( .A(\result_address[3][0] ), .B(remove_enable[3]), .C(
        \result_address[3][3] ), .Y(n273) );
  NAND3X1 U265 ( .A(\result_address[5][0] ), .B(remove_enable[5]), .C(
        \result_address[5][3] ), .Y(n151) );
  OAI21X1 U266 ( .A(n158), .B(n221), .C(n274), .Y(n269) );
  AOI22X1 U267 ( .A(n223), .B(n161), .C(n224), .D(n163), .Y(n274) );
  INVX1 U268 ( .A(n275), .Y(n163) );
  NAND3X1 U269 ( .A(\result_address[1][0] ), .B(remove_enable[1]), .C(
        \result_address[1][3] ), .Y(n275) );
  INVX1 U270 ( .A(n276), .Y(n161) );
  NAND3X1 U271 ( .A(\result_address[0][0] ), .B(remove_enable[0]), .C(
        \result_address[0][3] ), .Y(n276) );
  NAND3X1 U272 ( .A(\result_address[2][0] ), .B(remove_enable[2]), .C(
        \result_address[2][3] ), .Y(n158) );
  OR2X1 U273 ( .A(n277), .B(n278), .Y(dependency_remove[10]) );
  OAI21X1 U274 ( .A(n167), .B(n217), .C(n279), .Y(n278) );
  AOI22X1 U275 ( .A(n219), .B(n169), .C(n220), .D(n170), .Y(n279) );
  INVX1 U276 ( .A(n280), .Y(n170) );
  NAND3X1 U277 ( .A(remove_enable[4]), .B(n281), .C(\result_address[4][3] ), 
        .Y(n280) );
  NOR2X1 U278 ( .A(n251), .B(\result_address[4][2] ), .Y(n220) );
  INVX1 U279 ( .A(\result_address[4][1] ), .Y(n251) );
  INVX1 U280 ( .A(n282), .Y(n169) );
  NAND3X1 U281 ( .A(remove_enable[3]), .B(n283), .C(\result_address[3][3] ), 
        .Y(n282) );
  NOR2X1 U282 ( .A(n253), .B(\result_address[3][2] ), .Y(n219) );
  INVX1 U283 ( .A(\result_address[3][1] ), .Y(n253) );
  NAND2X1 U284 ( .A(\result_address[5][1] ), .B(n284), .Y(n217) );
  NAND3X1 U285 ( .A(remove_enable[5]), .B(n285), .C(\result_address[5][3] ), 
        .Y(n167) );
  OAI21X1 U286 ( .A(n171), .B(n221), .C(n286), .Y(n277) );
  AOI22X1 U287 ( .A(n223), .B(n173), .C(n224), .D(n174), .Y(n286) );
  INVX1 U288 ( .A(n287), .Y(n174) );
  NAND3X1 U289 ( .A(remove_enable[1]), .B(n288), .C(\result_address[1][3] ), 
        .Y(n287) );
  NOR2X1 U290 ( .A(n256), .B(\result_address[1][2] ), .Y(n224) );
  INVX1 U291 ( .A(\result_address[1][1] ), .Y(n256) );
  INVX1 U292 ( .A(n289), .Y(n173) );
  NAND3X1 U293 ( .A(remove_enable[0]), .B(n290), .C(\result_address[0][3] ), 
        .Y(n289) );
  NOR2X1 U294 ( .A(n258), .B(\result_address[0][2] ), .Y(n223) );
  INVX1 U295 ( .A(\result_address[0][1] ), .Y(n258) );
  NAND2X1 U296 ( .A(\result_address[2][1] ), .B(n291), .Y(n221) );
  NAND3X1 U297 ( .A(remove_enable[2]), .B(n292), .C(\result_address[2][3] ), 
        .Y(n171) );
  OR2X1 U298 ( .A(n293), .B(n294), .Y(dependency_remove[0]) );
  OAI21X1 U299 ( .A(n152), .B(n193), .C(n295), .Y(n294) );
  AOI22X1 U300 ( .A(n195), .B(n155), .C(n196), .D(n157), .Y(n295) );
  NOR2X1 U301 ( .A(\result_address[4][1] ), .B(\result_address[4][2] ), .Y(
        n157) );
  INVX1 U302 ( .A(n296), .Y(n196) );
  NAND3X1 U303 ( .A(n281), .B(n233), .C(remove_enable[4]), .Y(n296) );
  INVX1 U304 ( .A(\result_address[4][3] ), .Y(n233) );
  INVX1 U305 ( .A(\result_address[4][0] ), .Y(n281) );
  NOR2X1 U306 ( .A(\result_address[3][1] ), .B(\result_address[3][2] ), .Y(
        n155) );
  INVX1 U307 ( .A(n297), .Y(n195) );
  NAND3X1 U308 ( .A(n283), .B(n235), .C(remove_enable[3]), .Y(n297) );
  INVX1 U309 ( .A(\result_address[3][3] ), .Y(n235) );
  INVX1 U310 ( .A(\result_address[3][0] ), .Y(n283) );
  NAND3X1 U311 ( .A(n285), .B(n236), .C(remove_enable[5]), .Y(n193) );
  INVX1 U312 ( .A(\result_address[5][3] ), .Y(n236) );
  INVX1 U313 ( .A(\result_address[5][0] ), .Y(n285) );
  NAND2X1 U314 ( .A(n266), .B(n284), .Y(n152) );
  INVX1 U315 ( .A(\result_address[5][2] ), .Y(n284) );
  INVX1 U316 ( .A(\result_address[5][1] ), .Y(n266) );
  OAI21X1 U317 ( .A(n159), .B(n197), .C(n298), .Y(n293) );
  AOI22X1 U318 ( .A(n199), .B(n162), .C(n200), .D(n164), .Y(n298) );
  NOR2X1 U319 ( .A(\result_address[1][1] ), .B(\result_address[1][2] ), .Y(
        n164) );
  INVX1 U320 ( .A(n299), .Y(n200) );
  NAND3X1 U321 ( .A(n288), .B(n239), .C(remove_enable[1]), .Y(n299) );
  INVX1 U322 ( .A(\result_address[1][3] ), .Y(n239) );
  INVX1 U323 ( .A(\result_address[1][0] ), .Y(n288) );
  NOR2X1 U324 ( .A(\result_address[0][1] ), .B(\result_address[0][2] ), .Y(
        n162) );
  INVX1 U325 ( .A(n300), .Y(n199) );
  NAND3X1 U326 ( .A(n290), .B(n241), .C(remove_enable[0]), .Y(n300) );
  INVX1 U327 ( .A(\result_address[0][3] ), .Y(n241) );
  INVX1 U328 ( .A(\result_address[0][0] ), .Y(n290) );
  NAND3X1 U329 ( .A(n292), .B(n242), .C(remove_enable[2]), .Y(n197) );
  INVX1 U330 ( .A(\result_address[2][3] ), .Y(n242) );
  INVX1 U331 ( .A(\result_address[2][0] ), .Y(n292) );
  NAND2X1 U332 ( .A(n268), .B(n291), .Y(n159) );
  INVX1 U333 ( .A(\result_address[2][2] ), .Y(n291) );
  INVX1 U334 ( .A(\result_address[2][1] ), .Y(n268) );
endmodule

