
module upDownCounter_15 ( clk, n_rst, up, down, count_out );
  output [3:0] count_out;
  input clk, n_rst, up, down;
  wire   n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n5, n6, n7, n8, n9, n10;

  DFFSR \count_out_reg[0]  ( .D(n25), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[0]) );
  DFFSR \count_out_reg[1]  ( .D(n24), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[1]) );
  DFFSR \count_out_reg[2]  ( .D(n23), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[2]) );
  DFFSR \count_out_reg[3]  ( .D(n22), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[3]) );
  OAI22X1 U13 ( .A(n11), .B(n7), .C(n12), .D(n9), .Y(n22) );
  AOI22X1 U14 ( .A(n13), .B(n6), .C(count_out[3]), .D(n14), .Y(n11) );
  NAND3X1 U15 ( .A(up), .B(count_out[2]), .C(n5), .Y(n14) );
  NOR2X1 U16 ( .A(count_out[3]), .B(n8), .Y(n13) );
  OAI21X1 U17 ( .A(n16), .B(n17), .C(n18), .Y(n23) );
  OAI21X1 U18 ( .A(n15), .B(n19), .C(count_out[2]), .Y(n18) );
  NAND2X1 U19 ( .A(n12), .B(up), .Y(n19) );
  NAND2X1 U20 ( .A(count_out[1]), .B(count_out[0]), .Y(n15) );
  NAND2X1 U21 ( .A(n12), .B(n8), .Y(n17) );
  NAND3X1 U22 ( .A(count_out[1]), .B(count_out[0]), .C(up), .Y(n16) );
  XNOR2X1 U23 ( .A(count_out[1]), .B(n20), .Y(n24) );
  NAND3X1 U24 ( .A(n12), .B(count_out[0]), .C(up), .Y(n20) );
  XNOR2X1 U25 ( .A(count_out[0]), .B(n7), .Y(n25) );
  OAI21X1 U26 ( .A(down), .B(n10), .C(n21), .Y(n12) );
  NAND3X1 U27 ( .A(count_out[0]), .B(n10), .C(down), .Y(n21) );
  INVX2 U7 ( .A(n15), .Y(n5) );
  INVX2 U8 ( .A(n16), .Y(n6) );
  INVX2 U9 ( .A(n12), .Y(n7) );
  INVX2 U10 ( .A(count_out[2]), .Y(n8) );
  INVX2 U11 ( .A(count_out[3]), .Y(n9) );
  INVX2 U12 ( .A(up), .Y(n10) );
endmodule


module upDownCounter_14 ( clk, n_rst, up, down, count_out );
  output [3:0] count_out;
  input clk, n_rst, up, down;
  wire   n5, n6, n7, n8, n9, n10, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40;

  DFFSR \count_out_reg[0]  ( .D(n26), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[0]) );
  DFFSR \count_out_reg[1]  ( .D(n27), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[1]) );
  DFFSR \count_out_reg[2]  ( .D(n28), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[2]) );
  DFFSR \count_out_reg[3]  ( .D(n29), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[3]) );
  OAI22X1 U13 ( .A(n40), .B(n7), .C(n39), .D(n9), .Y(n29) );
  AOI22X1 U14 ( .A(n38), .B(n6), .C(count_out[3]), .D(n37), .Y(n40) );
  NAND3X1 U15 ( .A(up), .B(count_out[2]), .C(n5), .Y(n37) );
  NOR2X1 U16 ( .A(count_out[3]), .B(n8), .Y(n38) );
  OAI21X1 U17 ( .A(n35), .B(n34), .C(n33), .Y(n28) );
  OAI21X1 U18 ( .A(n36), .B(n32), .C(count_out[2]), .Y(n33) );
  NAND2X1 U19 ( .A(n39), .B(up), .Y(n32) );
  NAND2X1 U20 ( .A(count_out[1]), .B(count_out[0]), .Y(n36) );
  NAND2X1 U21 ( .A(n39), .B(n8), .Y(n34) );
  NAND3X1 U22 ( .A(count_out[1]), .B(count_out[0]), .C(up), .Y(n35) );
  XNOR2X1 U23 ( .A(count_out[1]), .B(n31), .Y(n27) );
  NAND3X1 U24 ( .A(n39), .B(count_out[0]), .C(up), .Y(n31) );
  XNOR2X1 U25 ( .A(count_out[0]), .B(n7), .Y(n26) );
  OAI21X1 U26 ( .A(down), .B(n10), .C(n30), .Y(n39) );
  NAND3X1 U27 ( .A(count_out[0]), .B(n10), .C(down), .Y(n30) );
  INVX2 U7 ( .A(n36), .Y(n5) );
  INVX2 U8 ( .A(n35), .Y(n6) );
  INVX2 U9 ( .A(n39), .Y(n7) );
  INVX2 U10 ( .A(count_out[2]), .Y(n8) );
  INVX2 U11 ( .A(count_out[3]), .Y(n9) );
  INVX2 U12 ( .A(up), .Y(n10) );
endmodule


module upDownCounter_13 ( clk, n_rst, up, down, count_out );
  output [3:0] count_out;
  input clk, n_rst, up, down;
  wire   n5, n6, n7, n8, n9, n10, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40;

  DFFSR \count_out_reg[0]  ( .D(n26), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[0]) );
  DFFSR \count_out_reg[1]  ( .D(n27), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[1]) );
  DFFSR \count_out_reg[2]  ( .D(n28), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[2]) );
  DFFSR \count_out_reg[3]  ( .D(n29), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[3]) );
  OAI22X1 U13 ( .A(n40), .B(n7), .C(n39), .D(n9), .Y(n29) );
  AOI22X1 U14 ( .A(n38), .B(n6), .C(count_out[3]), .D(n37), .Y(n40) );
  NAND3X1 U15 ( .A(up), .B(count_out[2]), .C(n5), .Y(n37) );
  NOR2X1 U16 ( .A(count_out[3]), .B(n8), .Y(n38) );
  OAI21X1 U17 ( .A(n35), .B(n34), .C(n33), .Y(n28) );
  OAI21X1 U18 ( .A(n36), .B(n32), .C(count_out[2]), .Y(n33) );
  NAND2X1 U19 ( .A(n39), .B(up), .Y(n32) );
  NAND2X1 U20 ( .A(count_out[1]), .B(count_out[0]), .Y(n36) );
  NAND2X1 U21 ( .A(n39), .B(n8), .Y(n34) );
  NAND3X1 U22 ( .A(count_out[1]), .B(count_out[0]), .C(up), .Y(n35) );
  XNOR2X1 U23 ( .A(count_out[1]), .B(n31), .Y(n27) );
  NAND3X1 U24 ( .A(n39), .B(count_out[0]), .C(up), .Y(n31) );
  XNOR2X1 U25 ( .A(count_out[0]), .B(n7), .Y(n26) );
  OAI21X1 U26 ( .A(down), .B(n10), .C(n30), .Y(n39) );
  NAND3X1 U27 ( .A(count_out[0]), .B(n10), .C(down), .Y(n30) );
  INVX2 U7 ( .A(n36), .Y(n5) );
  INVX2 U8 ( .A(n35), .Y(n6) );
  INVX2 U9 ( .A(n39), .Y(n7) );
  INVX2 U10 ( .A(count_out[2]), .Y(n8) );
  INVX2 U11 ( .A(count_out[3]), .Y(n9) );
  INVX2 U12 ( .A(up), .Y(n10) );
endmodule


module upDownCounter_12 ( clk, n_rst, up, down, count_out );
  output [3:0] count_out;
  input clk, n_rst, up, down;
  wire   n5, n6, n7, n8, n9, n10, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40;

  DFFSR \count_out_reg[0]  ( .D(n26), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[0]) );
  DFFSR \count_out_reg[1]  ( .D(n27), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[1]) );
  DFFSR \count_out_reg[2]  ( .D(n28), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[2]) );
  DFFSR \count_out_reg[3]  ( .D(n29), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[3]) );
  OAI22X1 U13 ( .A(n40), .B(n7), .C(n39), .D(n9), .Y(n29) );
  AOI22X1 U14 ( .A(n38), .B(n6), .C(count_out[3]), .D(n37), .Y(n40) );
  NAND3X1 U15 ( .A(up), .B(count_out[2]), .C(n5), .Y(n37) );
  NOR2X1 U16 ( .A(count_out[3]), .B(n8), .Y(n38) );
  OAI21X1 U17 ( .A(n35), .B(n34), .C(n33), .Y(n28) );
  OAI21X1 U18 ( .A(n36), .B(n32), .C(count_out[2]), .Y(n33) );
  NAND2X1 U19 ( .A(n39), .B(up), .Y(n32) );
  NAND2X1 U20 ( .A(count_out[1]), .B(count_out[0]), .Y(n36) );
  NAND2X1 U21 ( .A(n39), .B(n8), .Y(n34) );
  NAND3X1 U22 ( .A(count_out[1]), .B(count_out[0]), .C(up), .Y(n35) );
  XNOR2X1 U23 ( .A(count_out[1]), .B(n31), .Y(n27) );
  NAND3X1 U24 ( .A(n39), .B(count_out[0]), .C(up), .Y(n31) );
  XNOR2X1 U25 ( .A(count_out[0]), .B(n7), .Y(n26) );
  OAI21X1 U26 ( .A(down), .B(n10), .C(n30), .Y(n39) );
  NAND3X1 U27 ( .A(count_out[0]), .B(n10), .C(down), .Y(n30) );
  INVX2 U7 ( .A(n36), .Y(n5) );
  INVX2 U8 ( .A(n35), .Y(n6) );
  INVX2 U9 ( .A(n39), .Y(n7) );
  INVX2 U10 ( .A(count_out[2]), .Y(n8) );
  INVX2 U11 ( .A(count_out[3]), .Y(n9) );
  INVX2 U12 ( .A(up), .Y(n10) );
endmodule


module upDownCounter_11 ( clk, n_rst, up, down, count_out );
  output [3:0] count_out;
  input clk, n_rst, up, down;
  wire   n5, n6, n7, n8, n9, n10, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40;

  DFFSR \count_out_reg[0]  ( .D(n26), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[0]) );
  DFFSR \count_out_reg[1]  ( .D(n27), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[1]) );
  DFFSR \count_out_reg[2]  ( .D(n28), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[2]) );
  DFFSR \count_out_reg[3]  ( .D(n29), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[3]) );
  OAI22X1 U13 ( .A(n40), .B(n7), .C(n39), .D(n9), .Y(n29) );
  AOI22X1 U14 ( .A(n38), .B(n6), .C(count_out[3]), .D(n37), .Y(n40) );
  NAND3X1 U15 ( .A(up), .B(count_out[2]), .C(n5), .Y(n37) );
  NOR2X1 U16 ( .A(count_out[3]), .B(n8), .Y(n38) );
  OAI21X1 U17 ( .A(n35), .B(n34), .C(n33), .Y(n28) );
  OAI21X1 U18 ( .A(n36), .B(n32), .C(count_out[2]), .Y(n33) );
  NAND2X1 U19 ( .A(n39), .B(up), .Y(n32) );
  NAND2X1 U20 ( .A(count_out[1]), .B(count_out[0]), .Y(n36) );
  NAND2X1 U21 ( .A(n39), .B(n8), .Y(n34) );
  NAND3X1 U22 ( .A(count_out[1]), .B(count_out[0]), .C(up), .Y(n35) );
  XNOR2X1 U23 ( .A(count_out[1]), .B(n31), .Y(n27) );
  NAND3X1 U24 ( .A(n39), .B(count_out[0]), .C(up), .Y(n31) );
  XNOR2X1 U25 ( .A(count_out[0]), .B(n7), .Y(n26) );
  OAI21X1 U26 ( .A(down), .B(n10), .C(n30), .Y(n39) );
  NAND3X1 U27 ( .A(count_out[0]), .B(n10), .C(down), .Y(n30) );
  INVX2 U7 ( .A(n36), .Y(n5) );
  INVX2 U8 ( .A(n35), .Y(n6) );
  INVX2 U9 ( .A(n39), .Y(n7) );
  INVX2 U10 ( .A(count_out[2]), .Y(n8) );
  INVX2 U11 ( .A(count_out[3]), .Y(n9) );
  INVX2 U12 ( .A(up), .Y(n10) );
endmodule


module upDownCounter_10 ( clk, n_rst, up, down, count_out );
  output [3:0] count_out;
  input clk, n_rst, up, down;
  wire   n5, n6, n7, n8, n9, n10, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40;

  DFFSR \count_out_reg[0]  ( .D(n26), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[0]) );
  DFFSR \count_out_reg[1]  ( .D(n27), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[1]) );
  DFFSR \count_out_reg[2]  ( .D(n28), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[2]) );
  DFFSR \count_out_reg[3]  ( .D(n29), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[3]) );
  OAI22X1 U13 ( .A(n40), .B(n7), .C(n39), .D(n9), .Y(n29) );
  AOI22X1 U14 ( .A(n38), .B(n6), .C(count_out[3]), .D(n37), .Y(n40) );
  NAND3X1 U15 ( .A(up), .B(count_out[2]), .C(n5), .Y(n37) );
  NOR2X1 U16 ( .A(count_out[3]), .B(n8), .Y(n38) );
  OAI21X1 U17 ( .A(n35), .B(n34), .C(n33), .Y(n28) );
  OAI21X1 U18 ( .A(n36), .B(n32), .C(count_out[2]), .Y(n33) );
  NAND2X1 U19 ( .A(n39), .B(up), .Y(n32) );
  NAND2X1 U20 ( .A(count_out[1]), .B(count_out[0]), .Y(n36) );
  NAND2X1 U21 ( .A(n39), .B(n8), .Y(n34) );
  NAND3X1 U22 ( .A(count_out[1]), .B(count_out[0]), .C(up), .Y(n35) );
  XNOR2X1 U23 ( .A(count_out[1]), .B(n31), .Y(n27) );
  NAND3X1 U24 ( .A(n39), .B(count_out[0]), .C(up), .Y(n31) );
  XNOR2X1 U25 ( .A(count_out[0]), .B(n7), .Y(n26) );
  OAI21X1 U26 ( .A(down), .B(n10), .C(n30), .Y(n39) );
  NAND3X1 U27 ( .A(count_out[0]), .B(n10), .C(down), .Y(n30) );
  INVX2 U7 ( .A(n36), .Y(n5) );
  INVX2 U8 ( .A(n35), .Y(n6) );
  INVX2 U9 ( .A(n39), .Y(n7) );
  INVX2 U10 ( .A(count_out[2]), .Y(n8) );
  INVX2 U11 ( .A(count_out[3]), .Y(n9) );
  INVX2 U12 ( .A(up), .Y(n10) );
endmodule


module upDownCounter_9 ( clk, n_rst, up, down, count_out );
  output [3:0] count_out;
  input clk, n_rst, up, down;
  wire   n5, n6, n7, n8, n9, n10, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40;

  DFFSR \count_out_reg[0]  ( .D(n26), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[0]) );
  DFFSR \count_out_reg[1]  ( .D(n27), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[1]) );
  DFFSR \count_out_reg[2]  ( .D(n28), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[2]) );
  DFFSR \count_out_reg[3]  ( .D(n29), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[3]) );
  OAI22X1 U13 ( .A(n40), .B(n7), .C(n39), .D(n9), .Y(n29) );
  AOI22X1 U14 ( .A(n38), .B(n6), .C(count_out[3]), .D(n37), .Y(n40) );
  NAND3X1 U15 ( .A(up), .B(count_out[2]), .C(n5), .Y(n37) );
  NOR2X1 U16 ( .A(count_out[3]), .B(n8), .Y(n38) );
  OAI21X1 U17 ( .A(n35), .B(n34), .C(n33), .Y(n28) );
  OAI21X1 U18 ( .A(n36), .B(n32), .C(count_out[2]), .Y(n33) );
  NAND2X1 U19 ( .A(n39), .B(up), .Y(n32) );
  NAND2X1 U20 ( .A(count_out[1]), .B(count_out[0]), .Y(n36) );
  NAND2X1 U21 ( .A(n39), .B(n8), .Y(n34) );
  NAND3X1 U22 ( .A(count_out[1]), .B(count_out[0]), .C(up), .Y(n35) );
  XNOR2X1 U23 ( .A(count_out[1]), .B(n31), .Y(n27) );
  NAND3X1 U24 ( .A(n39), .B(count_out[0]), .C(up), .Y(n31) );
  XNOR2X1 U25 ( .A(count_out[0]), .B(n7), .Y(n26) );
  OAI21X1 U26 ( .A(down), .B(n10), .C(n30), .Y(n39) );
  NAND3X1 U27 ( .A(count_out[0]), .B(n10), .C(down), .Y(n30) );
  INVX2 U7 ( .A(n36), .Y(n5) );
  INVX2 U8 ( .A(n35), .Y(n6) );
  INVX2 U9 ( .A(n39), .Y(n7) );
  INVX2 U10 ( .A(count_out[2]), .Y(n8) );
  INVX2 U11 ( .A(count_out[3]), .Y(n9) );
  INVX2 U12 ( .A(up), .Y(n10) );
endmodule


module upDownCounter_8 ( clk, n_rst, up, down, count_out );
  output [3:0] count_out;
  input clk, n_rst, up, down;
  wire   n5, n6, n7, n8, n9, n10, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40;

  DFFSR \count_out_reg[0]  ( .D(n26), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[0]) );
  DFFSR \count_out_reg[1]  ( .D(n27), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[1]) );
  DFFSR \count_out_reg[2]  ( .D(n28), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[2]) );
  DFFSR \count_out_reg[3]  ( .D(n29), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[3]) );
  OAI22X1 U13 ( .A(n40), .B(n7), .C(n39), .D(n9), .Y(n29) );
  AOI22X1 U14 ( .A(n38), .B(n6), .C(count_out[3]), .D(n37), .Y(n40) );
  NAND3X1 U15 ( .A(up), .B(count_out[2]), .C(n5), .Y(n37) );
  NOR2X1 U16 ( .A(count_out[3]), .B(n8), .Y(n38) );
  OAI21X1 U17 ( .A(n35), .B(n34), .C(n33), .Y(n28) );
  OAI21X1 U18 ( .A(n36), .B(n32), .C(count_out[2]), .Y(n33) );
  NAND2X1 U19 ( .A(n39), .B(up), .Y(n32) );
  NAND2X1 U20 ( .A(count_out[1]), .B(count_out[0]), .Y(n36) );
  NAND2X1 U21 ( .A(n39), .B(n8), .Y(n34) );
  NAND3X1 U22 ( .A(count_out[1]), .B(count_out[0]), .C(up), .Y(n35) );
  XNOR2X1 U23 ( .A(count_out[1]), .B(n31), .Y(n27) );
  NAND3X1 U24 ( .A(n39), .B(count_out[0]), .C(up), .Y(n31) );
  XNOR2X1 U25 ( .A(count_out[0]), .B(n7), .Y(n26) );
  OAI21X1 U26 ( .A(down), .B(n10), .C(n30), .Y(n39) );
  NAND3X1 U27 ( .A(count_out[0]), .B(n10), .C(down), .Y(n30) );
  INVX2 U7 ( .A(n36), .Y(n5) );
  INVX2 U8 ( .A(n35), .Y(n6) );
  INVX2 U9 ( .A(n39), .Y(n7) );
  INVX2 U10 ( .A(count_out[2]), .Y(n8) );
  INVX2 U11 ( .A(count_out[3]), .Y(n9) );
  INVX2 U12 ( .A(up), .Y(n10) );
endmodule


module upDownCounter_7 ( clk, n_rst, up, down, count_out );
  output [3:0] count_out;
  input clk, n_rst, up, down;
  wire   n5, n6, n7, n8, n9, n10, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40;

  DFFSR \count_out_reg[0]  ( .D(n26), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[0]) );
  DFFSR \count_out_reg[1]  ( .D(n27), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[1]) );
  DFFSR \count_out_reg[2]  ( .D(n28), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[2]) );
  DFFSR \count_out_reg[3]  ( .D(n29), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[3]) );
  OAI22X1 U13 ( .A(n40), .B(n7), .C(n39), .D(n9), .Y(n29) );
  AOI22X1 U14 ( .A(n38), .B(n6), .C(count_out[3]), .D(n37), .Y(n40) );
  NAND3X1 U15 ( .A(up), .B(count_out[2]), .C(n5), .Y(n37) );
  NOR2X1 U16 ( .A(count_out[3]), .B(n8), .Y(n38) );
  OAI21X1 U17 ( .A(n35), .B(n34), .C(n33), .Y(n28) );
  OAI21X1 U18 ( .A(n36), .B(n32), .C(count_out[2]), .Y(n33) );
  NAND2X1 U19 ( .A(n39), .B(up), .Y(n32) );
  NAND2X1 U20 ( .A(count_out[1]), .B(count_out[0]), .Y(n36) );
  NAND2X1 U21 ( .A(n39), .B(n8), .Y(n34) );
  NAND3X1 U22 ( .A(count_out[1]), .B(count_out[0]), .C(up), .Y(n35) );
  XNOR2X1 U23 ( .A(count_out[1]), .B(n31), .Y(n27) );
  NAND3X1 U24 ( .A(n39), .B(count_out[0]), .C(up), .Y(n31) );
  XNOR2X1 U25 ( .A(count_out[0]), .B(n7), .Y(n26) );
  OAI21X1 U26 ( .A(down), .B(n10), .C(n30), .Y(n39) );
  NAND3X1 U27 ( .A(count_out[0]), .B(n10), .C(down), .Y(n30) );
  INVX2 U7 ( .A(n36), .Y(n5) );
  INVX2 U8 ( .A(n35), .Y(n6) );
  INVX2 U9 ( .A(n39), .Y(n7) );
  INVX2 U10 ( .A(count_out[2]), .Y(n8) );
  INVX2 U11 ( .A(count_out[3]), .Y(n9) );
  INVX2 U12 ( .A(up), .Y(n10) );
endmodule


module upDownCounter_6 ( clk, n_rst, up, down, count_out );
  output [3:0] count_out;
  input clk, n_rst, up, down;
  wire   n5, n6, n7, n8, n9, n10, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40;

  DFFSR \count_out_reg[0]  ( .D(n26), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[0]) );
  DFFSR \count_out_reg[1]  ( .D(n27), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[1]) );
  DFFSR \count_out_reg[2]  ( .D(n28), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[2]) );
  DFFSR \count_out_reg[3]  ( .D(n29), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[3]) );
  OAI22X1 U13 ( .A(n40), .B(n7), .C(n39), .D(n9), .Y(n29) );
  AOI22X1 U14 ( .A(n38), .B(n6), .C(count_out[3]), .D(n37), .Y(n40) );
  NAND3X1 U15 ( .A(up), .B(count_out[2]), .C(n5), .Y(n37) );
  NOR2X1 U16 ( .A(count_out[3]), .B(n8), .Y(n38) );
  OAI21X1 U17 ( .A(n35), .B(n34), .C(n33), .Y(n28) );
  OAI21X1 U18 ( .A(n36), .B(n32), .C(count_out[2]), .Y(n33) );
  NAND2X1 U19 ( .A(n39), .B(up), .Y(n32) );
  NAND2X1 U20 ( .A(count_out[1]), .B(count_out[0]), .Y(n36) );
  NAND2X1 U21 ( .A(n39), .B(n8), .Y(n34) );
  NAND3X1 U22 ( .A(count_out[1]), .B(count_out[0]), .C(up), .Y(n35) );
  XNOR2X1 U23 ( .A(count_out[1]), .B(n31), .Y(n27) );
  NAND3X1 U24 ( .A(n39), .B(count_out[0]), .C(up), .Y(n31) );
  XNOR2X1 U25 ( .A(count_out[0]), .B(n7), .Y(n26) );
  OAI21X1 U26 ( .A(down), .B(n10), .C(n30), .Y(n39) );
  NAND3X1 U27 ( .A(count_out[0]), .B(n10), .C(down), .Y(n30) );
  INVX2 U7 ( .A(n36), .Y(n5) );
  INVX2 U8 ( .A(n35), .Y(n6) );
  INVX2 U9 ( .A(n39), .Y(n7) );
  INVX2 U10 ( .A(count_out[2]), .Y(n8) );
  INVX2 U11 ( .A(count_out[3]), .Y(n9) );
  INVX2 U12 ( .A(up), .Y(n10) );
endmodule


module upDownCounter_5 ( clk, n_rst, up, down, count_out );
  output [3:0] count_out;
  input clk, n_rst, up, down;
  wire   n5, n6, n7, n8, n9, n10, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40;

  DFFSR \count_out_reg[0]  ( .D(n26), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[0]) );
  DFFSR \count_out_reg[1]  ( .D(n27), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[1]) );
  DFFSR \count_out_reg[2]  ( .D(n28), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[2]) );
  DFFSR \count_out_reg[3]  ( .D(n29), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[3]) );
  OAI22X1 U13 ( .A(n40), .B(n7), .C(n39), .D(n9), .Y(n29) );
  AOI22X1 U14 ( .A(n38), .B(n6), .C(count_out[3]), .D(n37), .Y(n40) );
  NAND3X1 U15 ( .A(up), .B(count_out[2]), .C(n5), .Y(n37) );
  NOR2X1 U16 ( .A(count_out[3]), .B(n8), .Y(n38) );
  OAI21X1 U17 ( .A(n35), .B(n34), .C(n33), .Y(n28) );
  OAI21X1 U18 ( .A(n36), .B(n32), .C(count_out[2]), .Y(n33) );
  NAND2X1 U19 ( .A(n39), .B(up), .Y(n32) );
  NAND2X1 U20 ( .A(count_out[1]), .B(count_out[0]), .Y(n36) );
  NAND2X1 U21 ( .A(n39), .B(n8), .Y(n34) );
  NAND3X1 U22 ( .A(count_out[1]), .B(count_out[0]), .C(up), .Y(n35) );
  XNOR2X1 U23 ( .A(count_out[1]), .B(n31), .Y(n27) );
  NAND3X1 U24 ( .A(n39), .B(count_out[0]), .C(up), .Y(n31) );
  XNOR2X1 U25 ( .A(count_out[0]), .B(n7), .Y(n26) );
  OAI21X1 U26 ( .A(down), .B(n10), .C(n30), .Y(n39) );
  NAND3X1 U27 ( .A(count_out[0]), .B(n10), .C(down), .Y(n30) );
  INVX2 U7 ( .A(n36), .Y(n5) );
  INVX2 U8 ( .A(n35), .Y(n6) );
  INVX2 U9 ( .A(n39), .Y(n7) );
  INVX2 U10 ( .A(count_out[2]), .Y(n8) );
  INVX2 U11 ( .A(count_out[3]), .Y(n9) );
  INVX2 U12 ( .A(up), .Y(n10) );
endmodule


module upDownCounter_4 ( clk, n_rst, up, down, count_out );
  output [3:0] count_out;
  input clk, n_rst, up, down;
  wire   n5, n6, n7, n8, n9, n10, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40;

  DFFSR \count_out_reg[0]  ( .D(n26), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[0]) );
  DFFSR \count_out_reg[1]  ( .D(n27), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[1]) );
  DFFSR \count_out_reg[2]  ( .D(n28), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[2]) );
  DFFSR \count_out_reg[3]  ( .D(n29), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[3]) );
  OAI22X1 U13 ( .A(n40), .B(n7), .C(n39), .D(n9), .Y(n29) );
  AOI22X1 U14 ( .A(n38), .B(n6), .C(count_out[3]), .D(n37), .Y(n40) );
  NAND3X1 U15 ( .A(up), .B(count_out[2]), .C(n5), .Y(n37) );
  NOR2X1 U16 ( .A(count_out[3]), .B(n8), .Y(n38) );
  OAI21X1 U17 ( .A(n35), .B(n34), .C(n33), .Y(n28) );
  OAI21X1 U18 ( .A(n36), .B(n32), .C(count_out[2]), .Y(n33) );
  NAND2X1 U19 ( .A(n39), .B(up), .Y(n32) );
  NAND2X1 U20 ( .A(count_out[1]), .B(count_out[0]), .Y(n36) );
  NAND2X1 U21 ( .A(n39), .B(n8), .Y(n34) );
  NAND3X1 U22 ( .A(count_out[1]), .B(count_out[0]), .C(up), .Y(n35) );
  XNOR2X1 U23 ( .A(count_out[1]), .B(n31), .Y(n27) );
  NAND3X1 U24 ( .A(n39), .B(count_out[0]), .C(up), .Y(n31) );
  XNOR2X1 U25 ( .A(count_out[0]), .B(n7), .Y(n26) );
  OAI21X1 U26 ( .A(down), .B(n10), .C(n30), .Y(n39) );
  NAND3X1 U27 ( .A(count_out[0]), .B(n10), .C(down), .Y(n30) );
  INVX2 U7 ( .A(n36), .Y(n5) );
  INVX2 U8 ( .A(n35), .Y(n6) );
  INVX2 U9 ( .A(n39), .Y(n7) );
  INVX2 U10 ( .A(count_out[2]), .Y(n8) );
  INVX2 U11 ( .A(count_out[3]), .Y(n9) );
  INVX2 U12 ( .A(up), .Y(n10) );
endmodule


module upDownCounter_3 ( clk, n_rst, up, down, count_out );
  output [3:0] count_out;
  input clk, n_rst, up, down;
  wire   n5, n6, n7, n8, n9, n10, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40;

  DFFSR \count_out_reg[0]  ( .D(n26), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[0]) );
  DFFSR \count_out_reg[1]  ( .D(n27), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[1]) );
  DFFSR \count_out_reg[2]  ( .D(n28), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[2]) );
  DFFSR \count_out_reg[3]  ( .D(n29), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[3]) );
  OAI22X1 U13 ( .A(n40), .B(n7), .C(n39), .D(n9), .Y(n29) );
  AOI22X1 U14 ( .A(n38), .B(n6), .C(count_out[3]), .D(n37), .Y(n40) );
  NAND3X1 U15 ( .A(up), .B(count_out[2]), .C(n5), .Y(n37) );
  NOR2X1 U16 ( .A(count_out[3]), .B(n8), .Y(n38) );
  OAI21X1 U17 ( .A(n35), .B(n34), .C(n33), .Y(n28) );
  OAI21X1 U18 ( .A(n36), .B(n32), .C(count_out[2]), .Y(n33) );
  NAND2X1 U19 ( .A(n39), .B(up), .Y(n32) );
  NAND2X1 U20 ( .A(count_out[1]), .B(count_out[0]), .Y(n36) );
  NAND2X1 U21 ( .A(n39), .B(n8), .Y(n34) );
  NAND3X1 U22 ( .A(count_out[1]), .B(count_out[0]), .C(up), .Y(n35) );
  XNOR2X1 U23 ( .A(count_out[1]), .B(n31), .Y(n27) );
  NAND3X1 U24 ( .A(n39), .B(count_out[0]), .C(up), .Y(n31) );
  XNOR2X1 U25 ( .A(count_out[0]), .B(n7), .Y(n26) );
  OAI21X1 U26 ( .A(down), .B(n10), .C(n30), .Y(n39) );
  NAND3X1 U27 ( .A(count_out[0]), .B(n10), .C(down), .Y(n30) );
  INVX2 U7 ( .A(n36), .Y(n5) );
  INVX2 U8 ( .A(n35), .Y(n6) );
  INVX2 U9 ( .A(n39), .Y(n7) );
  INVX2 U10 ( .A(count_out[2]), .Y(n8) );
  INVX2 U11 ( .A(count_out[3]), .Y(n9) );
  INVX2 U12 ( .A(up), .Y(n10) );
endmodule


module upDownCounter_2 ( clk, n_rst, up, down, count_out );
  output [3:0] count_out;
  input clk, n_rst, up, down;
  wire   n5, n6, n7, n8, n9, n10, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40;

  DFFSR \count_out_reg[0]  ( .D(n26), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[0]) );
  DFFSR \count_out_reg[1]  ( .D(n27), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[1]) );
  DFFSR \count_out_reg[2]  ( .D(n28), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[2]) );
  DFFSR \count_out_reg[3]  ( .D(n29), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[3]) );
  OAI22X1 U13 ( .A(n40), .B(n7), .C(n39), .D(n9), .Y(n29) );
  AOI22X1 U14 ( .A(n38), .B(n6), .C(count_out[3]), .D(n37), .Y(n40) );
  NAND3X1 U15 ( .A(up), .B(count_out[2]), .C(n5), .Y(n37) );
  NOR2X1 U16 ( .A(count_out[3]), .B(n8), .Y(n38) );
  OAI21X1 U17 ( .A(n35), .B(n34), .C(n33), .Y(n28) );
  OAI21X1 U18 ( .A(n36), .B(n32), .C(count_out[2]), .Y(n33) );
  NAND2X1 U19 ( .A(n39), .B(up), .Y(n32) );
  NAND2X1 U20 ( .A(count_out[1]), .B(count_out[0]), .Y(n36) );
  NAND2X1 U21 ( .A(n39), .B(n8), .Y(n34) );
  NAND3X1 U22 ( .A(count_out[1]), .B(count_out[0]), .C(up), .Y(n35) );
  XNOR2X1 U23 ( .A(count_out[1]), .B(n31), .Y(n27) );
  NAND3X1 U24 ( .A(n39), .B(count_out[0]), .C(up), .Y(n31) );
  XNOR2X1 U25 ( .A(count_out[0]), .B(n7), .Y(n26) );
  OAI21X1 U26 ( .A(down), .B(n10), .C(n30), .Y(n39) );
  NAND3X1 U27 ( .A(count_out[0]), .B(n10), .C(down), .Y(n30) );
  INVX2 U7 ( .A(n36), .Y(n5) );
  INVX2 U8 ( .A(n35), .Y(n6) );
  INVX2 U9 ( .A(n39), .Y(n7) );
  INVX2 U10 ( .A(count_out[2]), .Y(n8) );
  INVX2 U11 ( .A(count_out[3]), .Y(n9) );
  INVX2 U12 ( .A(up), .Y(n10) );
endmodule


module upDownCounter_1 ( clk, n_rst, up, down, count_out );
  output [3:0] count_out;
  input clk, n_rst, up, down;
  wire   n5, n6, n7, n8, n9, n10, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40;

  DFFSR \count_out_reg[0]  ( .D(n26), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[0]) );
  DFFSR \count_out_reg[1]  ( .D(n27), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[1]) );
  DFFSR \count_out_reg[2]  ( .D(n28), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[2]) );
  DFFSR \count_out_reg[3]  ( .D(n29), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[3]) );
  OAI22X1 U13 ( .A(n40), .B(n7), .C(n39), .D(n9), .Y(n29) );
  AOI22X1 U14 ( .A(n38), .B(n6), .C(count_out[3]), .D(n37), .Y(n40) );
  NAND3X1 U15 ( .A(up), .B(count_out[2]), .C(n5), .Y(n37) );
  NOR2X1 U16 ( .A(count_out[3]), .B(n8), .Y(n38) );
  OAI21X1 U17 ( .A(n35), .B(n34), .C(n33), .Y(n28) );
  OAI21X1 U18 ( .A(n36), .B(n32), .C(count_out[2]), .Y(n33) );
  NAND2X1 U19 ( .A(n39), .B(up), .Y(n32) );
  NAND2X1 U20 ( .A(count_out[1]), .B(count_out[0]), .Y(n36) );
  NAND2X1 U21 ( .A(n39), .B(n8), .Y(n34) );
  NAND3X1 U22 ( .A(count_out[1]), .B(count_out[0]), .C(up), .Y(n35) );
  XNOR2X1 U23 ( .A(count_out[1]), .B(n31), .Y(n27) );
  NAND3X1 U24 ( .A(n39), .B(count_out[0]), .C(up), .Y(n31) );
  XNOR2X1 U25 ( .A(count_out[0]), .B(n7), .Y(n26) );
  OAI21X1 U26 ( .A(down), .B(n10), .C(n30), .Y(n39) );
  NAND3X1 U27 ( .A(count_out[0]), .B(n10), .C(down), .Y(n30) );
  INVX2 U7 ( .A(n36), .Y(n5) );
  INVX2 U8 ( .A(n35), .Y(n6) );
  INVX2 U9 ( .A(n39), .Y(n7) );
  INVX2 U10 ( .A(count_out[2]), .Y(n8) );
  INVX2 U11 ( .A(count_out[3]), .Y(n9) );
  INVX2 U12 ( .A(up), .Y(n10) );
endmodule


module upDownCounter_0 ( clk, n_rst, up, down, count_out );
  output [3:0] count_out;
  input clk, n_rst, up, down;
  wire   n5, n6, n7, n8, n9, n10, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40;

  DFFSR \count_out_reg[0]  ( .D(n26), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[0]) );
  DFFSR \count_out_reg[1]  ( .D(n27), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[1]) );
  DFFSR \count_out_reg[2]  ( .D(n28), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[2]) );
  DFFSR \count_out_reg[3]  ( .D(n29), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[3]) );
  OAI22X1 U13 ( .A(n40), .B(n7), .C(n39), .D(n9), .Y(n29) );
  AOI22X1 U14 ( .A(n38), .B(n6), .C(count_out[3]), .D(n37), .Y(n40) );
  NAND3X1 U15 ( .A(up), .B(count_out[2]), .C(n5), .Y(n37) );
  NOR2X1 U16 ( .A(count_out[3]), .B(n8), .Y(n38) );
  OAI21X1 U17 ( .A(n35), .B(n34), .C(n33), .Y(n28) );
  OAI21X1 U18 ( .A(n36), .B(n32), .C(count_out[2]), .Y(n33) );
  NAND2X1 U19 ( .A(n39), .B(up), .Y(n32) );
  NAND2X1 U20 ( .A(count_out[1]), .B(count_out[0]), .Y(n36) );
  NAND2X1 U21 ( .A(n39), .B(n8), .Y(n34) );
  NAND3X1 U22 ( .A(count_out[1]), .B(count_out[0]), .C(up), .Y(n35) );
  XNOR2X1 U23 ( .A(count_out[1]), .B(n31), .Y(n27) );
  NAND3X1 U24 ( .A(n39), .B(count_out[0]), .C(up), .Y(n31) );
  XNOR2X1 U25 ( .A(count_out[0]), .B(n7), .Y(n26) );
  OAI21X1 U26 ( .A(down), .B(n10), .C(n30), .Y(n39) );
  NAND3X1 U27 ( .A(count_out[0]), .B(n10), .C(down), .Y(n30) );
  INVX2 U7 ( .A(n36), .Y(n5) );
  INVX2 U8 ( .A(n35), .Y(n6) );
  INVX2 U9 ( .A(n39), .Y(n7) );
  INVX2 U10 ( .A(count_out[2]), .Y(n8) );
  INVX2 U11 ( .A(count_out[3]), .Y(n9) );
  INVX2 U12 ( .A(up), .Y(n10) );
endmodule


module flex_indexer_NUM_CNT_BITS2_1 ( clk, n_rst, clear, count_enable, 
        rollover_val, count_out, rollover_flag );
  input [1:0] rollover_val;
  output [1:0] count_out;
  input clk, n_rst, clear, count_enable;
  output rollover_flag;
  wire   n17, net4848, net5206, net5843, n1, n2, n3, n4, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16;
  wire   [1:0] nxt_count;
  assign rollover_flag = 1'b0;
  assign count_out[0] = net5843;

  DFFSR \count_out_reg[0]  ( .D(nxt_count[0]), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(n17) );
  DFFSR \count_out_reg[1]  ( .D(nxt_count[1]), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(count_out[1]) );
  INVX2 U6 ( .A(n1), .Y(n2) );
  BUFX4 U7 ( .A(n17), .Y(net5843) );
  INVX1 U8 ( .A(net5843), .Y(net4848) );
  AND2X1 U9 ( .A(n16), .B(n15), .Y(nxt_count[0]) );
  INVX1 U10 ( .A(net4848), .Y(net5206) );
  INVX1 U11 ( .A(count_out[1]), .Y(n1) );
  NAND2X1 U12 ( .A(n2), .B(count_enable), .Y(n3) );
  INVX2 U13 ( .A(clear), .Y(n15) );
  OAI21X1 U14 ( .A(n3), .B(net4848), .C(n15), .Y(n12) );
  INVX2 U15 ( .A(rollover_val[1]), .Y(n7) );
  XOR2X1 U16 ( .A(net4848), .B(rollover_val[0]), .Y(n4) );
  OAI21X1 U17 ( .A(n2), .B(n7), .C(n4), .Y(n8) );
  AOI22X1 U18 ( .A(n8), .B(count_enable), .C(n2), .D(n7), .Y(n9) );
  OAI21X1 U19 ( .A(count_enable), .B(n1), .C(n9), .Y(n10) );
  OAI21X1 U20 ( .A(n2), .B(net5206), .C(n10), .Y(n11) );
  NOR2X1 U21 ( .A(n12), .B(n11), .Y(nxt_count[1]) );
  XOR2X1 U22 ( .A(rollover_val[1]), .B(n2), .Y(n13) );
  OAI21X1 U23 ( .A(rollover_val[0]), .B(n13), .C(net4848), .Y(n14) );
  MUX2X1 U24 ( .B(net4848), .A(n14), .S(count_enable), .Y(n16) );
endmodule


module flex_indexer_NUM_CNT_BITS2_0 ( clk, n_rst, clear, count_enable, 
        rollover_val, count_out, rollover_flag );
  input [1:0] rollover_val;
  output [1:0] count_out;
  input clk, n_rst, clear, count_enable;
  output rollover_flag;
  wire   n26, n27, n1, n3, n4, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23;
  wire   [1:0] nxt_count;
  assign rollover_flag = 1'b0;

  DFFSR \count_out_reg[0]  ( .D(nxt_count[0]), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(n27) );
  DFFSR \count_out_reg[1]  ( .D(nxt_count[1]), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(n26) );
  INVX2 U6 ( .A(count_out[0]), .Y(n3) );
  INVX4 U7 ( .A(n8), .Y(count_out[0]) );
  INVX1 U8 ( .A(n19), .Y(nxt_count[1]) );
  INVX2 U9 ( .A(n4), .Y(n1) );
  BUFX4 U10 ( .A(n26), .Y(count_out[1]) );
  INVX1 U11 ( .A(n26), .Y(n4) );
  INVX2 U12 ( .A(n27), .Y(n8) );
  AND2X1 U13 ( .A(n23), .B(n22), .Y(nxt_count[0]) );
  INVX2 U14 ( .A(rollover_val[1]), .Y(n12) );
  XOR2X1 U15 ( .A(n3), .B(rollover_val[0]), .Y(n10) );
  NAND2X1 U16 ( .A(rollover_val[1]), .B(n4), .Y(n9) );
  NAND2X1 U17 ( .A(n10), .B(n9), .Y(n11) );
  AOI22X1 U18 ( .A(n1), .B(n12), .C(count_enable), .D(n11), .Y(n15) );
  NAND2X1 U19 ( .A(n1), .B(count_enable), .Y(n13) );
  NAND2X1 U20 ( .A(n15), .B(n14), .Y(n18) );
  INVX2 U21 ( .A(n13), .Y(n14) );
  AOI21X1 U22 ( .A(count_out[0]), .B(n14), .C(clear), .Y(n17) );
  OAI21X1 U23 ( .A(n15), .B(n3), .C(n4), .Y(n16) );
  NAND3X1 U24 ( .A(n18), .B(n17), .C(n16), .Y(n19) );
  XOR2X1 U25 ( .A(rollover_val[1]), .B(n1), .Y(n20) );
  OAI21X1 U26 ( .A(rollover_val[0]), .B(n20), .C(n3), .Y(n21) );
  MUX2X1 U27 ( .B(n3), .A(n21), .S(count_enable), .Y(n23) );
  INVX2 U28 ( .A(clear), .Y(n22) );
endmodule


module flex_fifo_WIDTH32_DEPTH4_BITS_WIDTH5_BITS_DEPTH2 ( clk, n_rst, r_enable, 
        w_enable, w_data, r_data, full, empty );
  input [31:0] w_data;
  output [31:0] r_data;
  input clk, n_rst, r_enable, w_enable;
  output full, empty;
  wire   N4, N5, _2_net_, \data[3][31] , \data[3][30] , \data[3][29] ,
         \data[3][28] , \data[3][27] , \data[3][26] , \data[3][25] ,
         \data[3][24] , \data[3][23] , \data[3][22] , \data[3][21] ,
         \data[3][20] , \data[3][19] , \data[3][18] , \data[3][17] ,
         \data[3][16] , \data[3][15] , \data[3][14] , \data[3][13] ,
         \data[3][12] , \data[3][11] , \data[3][10] , \data[3][9] ,
         \data[3][8] , \data[3][7] , \data[3][6] , \data[3][5] , \data[3][4] ,
         \data[3][3] , \data[3][2] , \data[3][1] , \data[3][0] , \data[2][31] ,
         \data[2][30] , \data[2][29] , \data[2][28] , \data[2][27] ,
         \data[2][26] , \data[2][25] , \data[2][24] , \data[2][23] ,
         \data[2][22] , \data[2][21] , \data[2][20] , \data[2][19] ,
         \data[2][18] , \data[2][17] , \data[2][16] , \data[2][15] ,
         \data[2][14] , \data[2][13] , \data[2][12] , \data[2][11] ,
         \data[2][10] , \data[2][9] , \data[2][8] , \data[2][7] , \data[2][6] ,
         \data[2][5] , \data[2][4] , \data[2][3] , \data[2][2] , \data[2][1] ,
         \data[2][0] , \data[1][31] , \data[1][30] , \data[1][29] ,
         \data[1][28] , \data[1][27] , \data[1][26] , \data[1][25] ,
         \data[1][24] , \data[1][23] , \data[1][22] , \data[1][21] ,
         \data[1][20] , \data[1][19] , \data[1][18] , \data[1][17] ,
         \data[1][16] , \data[1][15] , \data[1][14] , \data[1][13] ,
         \data[1][12] , \data[1][11] , \data[1][10] , \data[1][9] ,
         \data[1][8] , \data[1][7] , \data[1][6] , \data[1][5] , \data[1][4] ,
         \data[1][3] , \data[1][2] , \data[1][1] , \data[1][0] , \data[0][31] ,
         \data[0][30] , \data[0][29] , \data[0][28] , \data[0][27] ,
         \data[0][26] , \data[0][25] , \data[0][24] , \data[0][23] ,
         \data[0][22] , \data[0][21] , \data[0][20] , \data[0][19] ,
         \data[0][18] , \data[0][17] , \data[0][16] , \data[0][15] ,
         \data[0][14] , \data[0][13] , \data[0][12] , \data[0][11] ,
         \data[0][10] , \data[0][9] , \data[0][8] , \data[0][7] , \data[0][6] ,
         \data[0][5] , \data[0][4] , \data[0][3] , \data[0][2] , \data[0][1] ,
         \data[0][0] , \nxt_data[3][31] , \nxt_data[3][30] , \nxt_data[3][29] ,
         \nxt_data[3][28] , \nxt_data[3][27] , \nxt_data[3][26] ,
         \nxt_data[3][25] , \nxt_data[3][24] , \nxt_data[3][23] ,
         \nxt_data[3][22] , \nxt_data[3][21] , \nxt_data[3][20] ,
         \nxt_data[3][19] , \nxt_data[3][18] , \nxt_data[3][17] ,
         \nxt_data[3][16] , \nxt_data[3][15] , \nxt_data[3][14] ,
         \nxt_data[3][13] , \nxt_data[3][12] , \nxt_data[3][11] ,
         \nxt_data[3][10] , \nxt_data[3][9] , \nxt_data[3][8] ,
         \nxt_data[3][7] , \nxt_data[3][6] , \nxt_data[3][5] ,
         \nxt_data[3][4] , \nxt_data[3][3] , \nxt_data[3][2] ,
         \nxt_data[3][1] , \nxt_data[3][0] , \nxt_data[2][31] ,
         \nxt_data[2][30] , \nxt_data[2][29] , \nxt_data[2][28] ,
         \nxt_data[2][27] , \nxt_data[2][26] , \nxt_data[2][25] ,
         \nxt_data[2][24] , \nxt_data[2][23] , \nxt_data[2][22] ,
         \nxt_data[2][21] , \nxt_data[2][20] , \nxt_data[2][19] ,
         \nxt_data[2][18] , \nxt_data[2][17] , \nxt_data[2][16] ,
         \nxt_data[2][15] , \nxt_data[2][14] , \nxt_data[2][13] ,
         \nxt_data[2][12] , \nxt_data[2][11] , \nxt_data[2][10] ,
         \nxt_data[2][9] , \nxt_data[2][8] , \nxt_data[2][7] ,
         \nxt_data[2][6] , \nxt_data[2][5] , \nxt_data[2][4] ,
         \nxt_data[2][3] , \nxt_data[2][2] , \nxt_data[2][1] ,
         \nxt_data[2][0] , \nxt_data[1][31] , \nxt_data[1][30] ,
         \nxt_data[1][29] , \nxt_data[1][28] , \nxt_data[1][27] ,
         \nxt_data[1][26] , \nxt_data[1][25] , \nxt_data[1][24] ,
         \nxt_data[1][23] , \nxt_data[1][22] , \nxt_data[1][21] ,
         \nxt_data[1][20] , \nxt_data[1][19] , \nxt_data[1][18] ,
         \nxt_data[1][17] , \nxt_data[1][16] , \nxt_data[1][15] ,
         \nxt_data[1][14] , \nxt_data[1][13] , \nxt_data[1][12] ,
         \nxt_data[1][11] , \nxt_data[1][10] , \nxt_data[1][9] ,
         \nxt_data[1][8] , \nxt_data[1][7] , \nxt_data[1][6] ,
         \nxt_data[1][5] , \nxt_data[1][4] , \nxt_data[1][3] ,
         \nxt_data[1][2] , \nxt_data[1][1] , \nxt_data[1][0] ,
         \nxt_data[0][31] , \nxt_data[0][30] , \nxt_data[0][29] ,
         \nxt_data[0][28] , \nxt_data[0][27] , \nxt_data[0][26] ,
         \nxt_data[0][25] , \nxt_data[0][24] , \nxt_data[0][23] ,
         \nxt_data[0][22] , \nxt_data[0][21] , \nxt_data[0][20] ,
         \nxt_data[0][19] , \nxt_data[0][18] , \nxt_data[0][17] ,
         \nxt_data[0][16] , \nxt_data[0][15] , \nxt_data[0][14] ,
         \nxt_data[0][13] , \nxt_data[0][12] , \nxt_data[0][11] ,
         \nxt_data[0][10] , \nxt_data[0][9] , \nxt_data[0][8] ,
         \nxt_data[0][7] , \nxt_data[0][6] , \nxt_data[0][5] ,
         \nxt_data[0][4] , \nxt_data[0][3] , \nxt_data[0][2] ,
         \nxt_data[0][1] , \nxt_data[0][0] , N14, net2542, net4924, net4928,
         net4929, net4965, net4999, net5000, net5036, net5037, net5079,
         net5101, net5099, net5123, net5121, net5129, net5127, net5158,
         net5160, net5180, net5186, net5185, net5191, net5196, \C447/net5087 ,
         \C447/net5091 , \C447/net5067 , \C447/net5069 , \C447/net5071 ,
         \C447/net5073 , \C447/net5075 , net5841, net5133, net5211, net5035,
         net5842, net5201, n1, n2, n3, n4, n5, n6, n7, n8, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387;
  wire   [1:0] w_pointer;
  assign empty = N14;
  assign full = net2542;

  DFFSR \data_reg[3][31]  ( .D(\nxt_data[3][31] ), .CLK(clk), .R(n215), .S(
        1'b1), .Q(\data[3][31] ) );
  DFFSR \data_reg[3][30]  ( .D(\nxt_data[3][30] ), .CLK(clk), .R(n215), .S(
        1'b1), .Q(\data[3][30] ) );
  DFFSR \data_reg[3][29]  ( .D(\nxt_data[3][29] ), .CLK(clk), .R(n215), .S(
        1'b1), .Q(\data[3][29] ) );
  DFFSR \data_reg[3][28]  ( .D(\nxt_data[3][28] ), .CLK(clk), .R(n215), .S(
        1'b1), .Q(\data[3][28] ) );
  DFFSR \data_reg[3][27]  ( .D(\nxt_data[3][27] ), .CLK(clk), .R(n215), .S(
        1'b1), .Q(\data[3][27] ) );
  DFFSR \data_reg[3][26]  ( .D(\nxt_data[3][26] ), .CLK(clk), .R(n215), .S(
        1'b1), .Q(\data[3][26] ) );
  DFFSR \data_reg[3][25]  ( .D(\nxt_data[3][25] ), .CLK(clk), .R(n215), .S(
        1'b1), .Q(\data[3][25] ) );
  DFFSR \data_reg[3][24]  ( .D(\nxt_data[3][24] ), .CLK(clk), .R(n215), .S(
        1'b1), .Q(\data[3][24] ) );
  DFFSR \data_reg[3][23]  ( .D(\nxt_data[3][23] ), .CLK(clk), .R(n215), .S(
        1'b1), .Q(\data[3][23] ) );
  DFFSR \data_reg[3][22]  ( .D(\nxt_data[3][22] ), .CLK(clk), .R(n215), .S(
        1'b1), .Q(\data[3][22] ) );
  DFFSR \data_reg[3][21]  ( .D(\nxt_data[3][21] ), .CLK(clk), .R(n215), .S(
        1'b1), .Q(\data[3][21] ) );
  DFFSR \data_reg[3][20]  ( .D(\nxt_data[3][20] ), .CLK(clk), .R(n215), .S(
        1'b1), .Q(\data[3][20] ) );
  DFFSR \data_reg[3][19]  ( .D(\nxt_data[3][19] ), .CLK(clk), .R(n214), .S(
        1'b1), .Q(\data[3][19] ) );
  DFFSR \data_reg[3][18]  ( .D(\nxt_data[3][18] ), .CLK(clk), .R(n214), .S(
        1'b1), .Q(\data[3][18] ) );
  DFFSR \data_reg[3][17]  ( .D(\nxt_data[3][17] ), .CLK(clk), .R(n214), .S(
        1'b1), .Q(\data[3][17] ) );
  DFFSR \data_reg[3][16]  ( .D(\nxt_data[3][16] ), .CLK(clk), .R(n214), .S(
        1'b1), .Q(\data[3][16] ) );
  DFFSR \data_reg[3][15]  ( .D(\nxt_data[3][15] ), .CLK(clk), .R(n214), .S(
        1'b1), .Q(\data[3][15] ) );
  DFFSR \data_reg[3][14]  ( .D(\nxt_data[3][14] ), .CLK(clk), .R(n214), .S(
        1'b1), .Q(\data[3][14] ) );
  DFFSR \data_reg[3][13]  ( .D(\nxt_data[3][13] ), .CLK(clk), .R(n214), .S(
        1'b1), .Q(\data[3][13] ) );
  DFFSR \data_reg[3][12]  ( .D(\nxt_data[3][12] ), .CLK(clk), .R(n214), .S(
        1'b1), .Q(\data[3][12] ) );
  DFFSR \data_reg[3][11]  ( .D(\nxt_data[3][11] ), .CLK(clk), .R(n214), .S(
        1'b1), .Q(\data[3][11] ) );
  DFFSR \data_reg[3][10]  ( .D(\nxt_data[3][10] ), .CLK(clk), .R(n214), .S(
        1'b1), .Q(\data[3][10] ) );
  DFFSR \data_reg[3][9]  ( .D(\nxt_data[3][9] ), .CLK(clk), .R(n214), .S(1'b1), 
        .Q(\data[3][9] ) );
  DFFSR \data_reg[3][8]  ( .D(\nxt_data[3][8] ), .CLK(clk), .R(n214), .S(1'b1), 
        .Q(\data[3][8] ) );
  DFFSR \data_reg[3][7]  ( .D(\nxt_data[3][7] ), .CLK(clk), .R(n214), .S(1'b1), 
        .Q(\data[3][7] ) );
  DFFSR \data_reg[3][6]  ( .D(\nxt_data[3][6] ), .CLK(clk), .R(n214), .S(1'b1), 
        .Q(\data[3][6] ) );
  DFFSR \data_reg[3][5]  ( .D(\nxt_data[3][5] ), .CLK(clk), .R(n214), .S(1'b1), 
        .Q(\data[3][5] ) );
  DFFSR \data_reg[3][4]  ( .D(\nxt_data[3][4] ), .CLK(clk), .R(n214), .S(1'b1), 
        .Q(\data[3][4] ) );
  DFFSR \data_reg[3][3]  ( .D(\nxt_data[3][3] ), .CLK(clk), .R(n214), .S(1'b1), 
        .Q(\data[3][3] ) );
  DFFSR \data_reg[3][2]  ( .D(\nxt_data[3][2] ), .CLK(clk), .R(n214), .S(1'b1), 
        .Q(\data[3][2] ) );
  DFFSR \data_reg[3][1]  ( .D(\nxt_data[3][1] ), .CLK(clk), .R(n214), .S(1'b1), 
        .Q(\data[3][1] ) );
  DFFSR \data_reg[3][0]  ( .D(\nxt_data[3][0] ), .CLK(clk), .R(n214), .S(1'b1), 
        .Q(\data[3][0] ) );
  DFFSR \data_reg[2][31]  ( .D(\nxt_data[2][31] ), .CLK(clk), .R(n214), .S(
        1'b1), .Q(\data[2][31] ) );
  DFFSR \data_reg[2][30]  ( .D(\nxt_data[2][30] ), .CLK(clk), .R(n214), .S(
        1'b1), .Q(\data[2][30] ) );
  DFFSR \data_reg[2][29]  ( .D(\nxt_data[2][29] ), .CLK(clk), .R(n214), .S(
        1'b1), .Q(\data[2][29] ) );
  DFFSR \data_reg[2][28]  ( .D(\nxt_data[2][28] ), .CLK(clk), .R(n214), .S(
        1'b1), .Q(\data[2][28] ) );
  DFFSR \data_reg[2][27]  ( .D(\nxt_data[2][27] ), .CLK(clk), .R(n213), .S(
        1'b1), .Q(\data[2][27] ) );
  DFFSR \data_reg[2][26]  ( .D(\nxt_data[2][26] ), .CLK(clk), .R(n213), .S(
        1'b1), .Q(\data[2][26] ) );
  DFFSR \data_reg[2][25]  ( .D(\nxt_data[2][25] ), .CLK(clk), .R(n213), .S(
        1'b1), .Q(\data[2][25] ) );
  DFFSR \data_reg[2][24]  ( .D(\nxt_data[2][24] ), .CLK(clk), .R(n213), .S(
        1'b1), .Q(\data[2][24] ) );
  DFFSR \data_reg[2][23]  ( .D(\nxt_data[2][23] ), .CLK(clk), .R(n213), .S(
        1'b1), .Q(\data[2][23] ) );
  DFFSR \data_reg[2][22]  ( .D(\nxt_data[2][22] ), .CLK(clk), .R(n213), .S(
        1'b1), .Q(\data[2][22] ) );
  DFFSR \data_reg[2][21]  ( .D(\nxt_data[2][21] ), .CLK(clk), .R(n213), .S(
        1'b1), .Q(\data[2][21] ) );
  DFFSR \data_reg[2][20]  ( .D(\nxt_data[2][20] ), .CLK(clk), .R(n213), .S(
        1'b1), .Q(\data[2][20] ) );
  DFFSR \data_reg[2][19]  ( .D(\nxt_data[2][19] ), .CLK(clk), .R(n213), .S(
        1'b1), .Q(\data[2][19] ) );
  DFFSR \data_reg[2][18]  ( .D(\nxt_data[2][18] ), .CLK(clk), .R(n213), .S(
        1'b1), .Q(\data[2][18] ) );
  DFFSR \data_reg[2][17]  ( .D(\nxt_data[2][17] ), .CLK(clk), .R(n213), .S(
        1'b1), .Q(\data[2][17] ) );
  DFFSR \data_reg[2][16]  ( .D(\nxt_data[2][16] ), .CLK(clk), .R(n213), .S(
        1'b1), .Q(\data[2][16] ) );
  DFFSR \data_reg[2][15]  ( .D(\nxt_data[2][15] ), .CLK(clk), .R(n213), .S(
        1'b1), .Q(\data[2][15] ) );
  DFFSR \data_reg[2][14]  ( .D(\nxt_data[2][14] ), .CLK(clk), .R(n213), .S(
        1'b1), .Q(\data[2][14] ) );
  DFFSR \data_reg[2][13]  ( .D(\nxt_data[2][13] ), .CLK(clk), .R(n213), .S(
        1'b1), .Q(\data[2][13] ) );
  DFFSR \data_reg[2][12]  ( .D(\nxt_data[2][12] ), .CLK(clk), .R(n213), .S(
        1'b1), .Q(\data[2][12] ) );
  DFFSR \data_reg[2][11]  ( .D(\nxt_data[2][11] ), .CLK(clk), .R(n213), .S(
        1'b1), .Q(\data[2][11] ) );
  DFFSR \data_reg[2][10]  ( .D(\nxt_data[2][10] ), .CLK(clk), .R(n213), .S(
        1'b1), .Q(\data[2][10] ) );
  DFFSR \data_reg[2][9]  ( .D(\nxt_data[2][9] ), .CLK(clk), .R(n213), .S(1'b1), 
        .Q(\data[2][9] ) );
  DFFSR \data_reg[2][8]  ( .D(\nxt_data[2][8] ), .CLK(clk), .R(n213), .S(1'b1), 
        .Q(\data[2][8] ) );
  DFFSR \data_reg[2][7]  ( .D(\nxt_data[2][7] ), .CLK(clk), .R(n213), .S(1'b1), 
        .Q(\data[2][7] ) );
  DFFSR \data_reg[2][6]  ( .D(\nxt_data[2][6] ), .CLK(clk), .R(n213), .S(1'b1), 
        .Q(\data[2][6] ) );
  DFFSR \data_reg[2][5]  ( .D(\nxt_data[2][5] ), .CLK(clk), .R(n213), .S(1'b1), 
        .Q(\data[2][5] ) );
  DFFSR \data_reg[2][4]  ( .D(\nxt_data[2][4] ), .CLK(clk), .R(n213), .S(1'b1), 
        .Q(\data[2][4] ) );
  DFFSR \data_reg[2][3]  ( .D(\nxt_data[2][3] ), .CLK(clk), .R(n212), .S(1'b1), 
        .Q(\data[2][3] ) );
  DFFSR \data_reg[2][2]  ( .D(\nxt_data[2][2] ), .CLK(clk), .R(n212), .S(1'b1), 
        .Q(\data[2][2] ) );
  DFFSR \data_reg[2][1]  ( .D(\nxt_data[2][1] ), .CLK(clk), .R(n212), .S(1'b1), 
        .Q(\data[2][1] ) );
  DFFSR \data_reg[2][0]  ( .D(\nxt_data[2][0] ), .CLK(clk), .R(n212), .S(1'b1), 
        .Q(\data[2][0] ) );
  DFFSR \data_reg[1][31]  ( .D(\nxt_data[1][31] ), .CLK(clk), .R(n212), .S(
        1'b1), .Q(\data[1][31] ) );
  DFFSR \data_reg[1][30]  ( .D(\nxt_data[1][30] ), .CLK(clk), .R(n212), .S(
        1'b1), .Q(\data[1][30] ) );
  DFFSR \data_reg[1][29]  ( .D(\nxt_data[1][29] ), .CLK(clk), .R(n212), .S(
        1'b1), .Q(\data[1][29] ) );
  DFFSR \data_reg[1][28]  ( .D(\nxt_data[1][28] ), .CLK(clk), .R(n212), .S(
        1'b1), .Q(\data[1][28] ) );
  DFFSR \data_reg[1][27]  ( .D(\nxt_data[1][27] ), .CLK(clk), .R(n212), .S(
        1'b1), .Q(\data[1][27] ) );
  DFFSR \data_reg[1][26]  ( .D(\nxt_data[1][26] ), .CLK(clk), .R(n212), .S(
        1'b1), .Q(\data[1][26] ) );
  DFFSR \data_reg[1][25]  ( .D(\nxt_data[1][25] ), .CLK(clk), .R(n212), .S(
        1'b1), .Q(\data[1][25] ) );
  DFFSR \data_reg[1][24]  ( .D(\nxt_data[1][24] ), .CLK(clk), .R(n212), .S(
        1'b1), .Q(\data[1][24] ) );
  DFFSR \data_reg[1][23]  ( .D(\nxt_data[1][23] ), .CLK(clk), .R(n212), .S(
        1'b1), .Q(\data[1][23] ) );
  DFFSR \data_reg[1][22]  ( .D(\nxt_data[1][22] ), .CLK(clk), .R(n212), .S(
        1'b1), .Q(\data[1][22] ) );
  DFFSR \data_reg[1][21]  ( .D(\nxt_data[1][21] ), .CLK(clk), .R(n212), .S(
        1'b1), .Q(\data[1][21] ) );
  DFFSR \data_reg[1][20]  ( .D(\nxt_data[1][20] ), .CLK(clk), .R(n212), .S(
        1'b1), .Q(\data[1][20] ) );
  DFFSR \data_reg[1][19]  ( .D(\nxt_data[1][19] ), .CLK(clk), .R(n212), .S(
        1'b1), .Q(\data[1][19] ) );
  DFFSR \data_reg[1][18]  ( .D(\nxt_data[1][18] ), .CLK(clk), .R(n212), .S(
        1'b1), .Q(\data[1][18] ) );
  DFFSR \data_reg[1][17]  ( .D(\nxt_data[1][17] ), .CLK(clk), .R(n212), .S(
        1'b1), .Q(\data[1][17] ) );
  DFFSR \data_reg[1][16]  ( .D(\nxt_data[1][16] ), .CLK(clk), .R(n212), .S(
        1'b1), .Q(\data[1][16] ) );
  DFFSR \data_reg[1][15]  ( .D(\nxt_data[1][15] ), .CLK(clk), .R(n212), .S(
        1'b1), .Q(\data[1][15] ) );
  DFFSR \data_reg[1][14]  ( .D(\nxt_data[1][14] ), .CLK(clk), .R(n212), .S(
        1'b1), .Q(\data[1][14] ) );
  DFFSR \data_reg[1][13]  ( .D(\nxt_data[1][13] ), .CLK(clk), .R(n212), .S(
        1'b1), .Q(\data[1][13] ) );
  DFFSR \data_reg[1][12]  ( .D(\nxt_data[1][12] ), .CLK(clk), .R(n212), .S(
        1'b1), .Q(\data[1][12] ) );
  DFFSR \data_reg[1][11]  ( .D(\nxt_data[1][11] ), .CLK(clk), .R(n211), .S(
        1'b1), .Q(\data[1][11] ) );
  DFFSR \data_reg[1][10]  ( .D(\nxt_data[1][10] ), .CLK(clk), .R(n211), .S(
        1'b1), .Q(\data[1][10] ) );
  DFFSR \data_reg[1][9]  ( .D(\nxt_data[1][9] ), .CLK(clk), .R(n211), .S(1'b1), 
        .Q(\data[1][9] ) );
  DFFSR \data_reg[1][8]  ( .D(\nxt_data[1][8] ), .CLK(clk), .R(n211), .S(1'b1), 
        .Q(\data[1][8] ) );
  DFFSR \data_reg[1][7]  ( .D(\nxt_data[1][7] ), .CLK(clk), .R(n211), .S(1'b1), 
        .Q(\data[1][7] ) );
  DFFSR \data_reg[1][6]  ( .D(\nxt_data[1][6] ), .CLK(clk), .R(n211), .S(1'b1), 
        .Q(\data[1][6] ) );
  DFFSR \data_reg[1][5]  ( .D(\nxt_data[1][5] ), .CLK(clk), .R(n211), .S(1'b1), 
        .Q(\data[1][5] ) );
  DFFSR \data_reg[1][4]  ( .D(\nxt_data[1][4] ), .CLK(clk), .R(n211), .S(1'b1), 
        .Q(\data[1][4] ) );
  DFFSR \data_reg[1][3]  ( .D(\nxt_data[1][3] ), .CLK(clk), .R(n211), .S(1'b1), 
        .Q(\data[1][3] ) );
  DFFSR \data_reg[1][2]  ( .D(\nxt_data[1][2] ), .CLK(clk), .R(n211), .S(1'b1), 
        .Q(\data[1][2] ) );
  DFFSR \data_reg[1][1]  ( .D(\nxt_data[1][1] ), .CLK(clk), .R(n211), .S(1'b1), 
        .Q(\data[1][1] ) );
  DFFSR \data_reg[1][0]  ( .D(\nxt_data[1][0] ), .CLK(clk), .R(n211), .S(1'b1), 
        .Q(\data[1][0] ) );
  DFFSR \data_reg[0][31]  ( .D(\nxt_data[0][31] ), .CLK(clk), .R(n211), .S(
        1'b1), .Q(\data[0][31] ) );
  DFFSR \data_reg[0][30]  ( .D(\nxt_data[0][30] ), .CLK(clk), .R(n211), .S(
        1'b1), .Q(\data[0][30] ) );
  DFFSR \data_reg[0][29]  ( .D(\nxt_data[0][29] ), .CLK(clk), .R(n211), .S(
        1'b1), .Q(\data[0][29] ) );
  DFFSR \data_reg[0][28]  ( .D(\nxt_data[0][28] ), .CLK(clk), .R(n211), .S(
        1'b1), .Q(\data[0][28] ) );
  DFFSR \data_reg[0][27]  ( .D(\nxt_data[0][27] ), .CLK(clk), .R(n211), .S(
        1'b1), .Q(\data[0][27] ) );
  DFFSR \data_reg[0][26]  ( .D(\nxt_data[0][26] ), .CLK(clk), .R(n211), .S(
        1'b1), .Q(\data[0][26] ) );
  DFFSR \data_reg[0][25]  ( .D(\nxt_data[0][25] ), .CLK(clk), .R(n211), .S(
        1'b1), .Q(\data[0][25] ) );
  DFFSR \data_reg[0][24]  ( .D(\nxt_data[0][24] ), .CLK(clk), .R(n211), .S(
        1'b1), .Q(\data[0][24] ) );
  DFFSR \data_reg[0][23]  ( .D(\nxt_data[0][23] ), .CLK(clk), .R(n211), .S(
        1'b1), .Q(\data[0][23] ) );
  DFFSR \data_reg[0][22]  ( .D(\nxt_data[0][22] ), .CLK(clk), .R(n211), .S(
        1'b1), .Q(\data[0][22] ) );
  DFFSR \data_reg[0][21]  ( .D(\nxt_data[0][21] ), .CLK(clk), .R(n211), .S(
        1'b1), .Q(\data[0][21] ) );
  DFFSR \data_reg[0][20]  ( .D(\nxt_data[0][20] ), .CLK(clk), .R(n211), .S(
        1'b1), .Q(\data[0][20] ) );
  DFFSR \data_reg[0][19]  ( .D(\nxt_data[0][19] ), .CLK(clk), .R(n210), .S(
        1'b1), .Q(\data[0][19] ) );
  DFFSR \data_reg[0][18]  ( .D(\nxt_data[0][18] ), .CLK(clk), .R(n210), .S(
        1'b1), .Q(\data[0][18] ) );
  DFFSR \data_reg[0][17]  ( .D(\nxt_data[0][17] ), .CLK(clk), .R(n210), .S(
        1'b1), .Q(\data[0][17] ) );
  DFFSR \data_reg[0][16]  ( .D(\nxt_data[0][16] ), .CLK(clk), .R(n210), .S(
        1'b1), .Q(\data[0][16] ) );
  DFFSR \data_reg[0][15]  ( .D(\nxt_data[0][15] ), .CLK(clk), .R(n210), .S(
        1'b1), .Q(\data[0][15] ) );
  DFFSR \data_reg[0][14]  ( .D(\nxt_data[0][14] ), .CLK(clk), .R(n210), .S(
        1'b1), .Q(\data[0][14] ) );
  DFFSR \data_reg[0][13]  ( .D(\nxt_data[0][13] ), .CLK(clk), .R(n210), .S(
        1'b1), .Q(\data[0][13] ) );
  DFFSR \data_reg[0][12]  ( .D(\nxt_data[0][12] ), .CLK(clk), .R(n210), .S(
        1'b1), .Q(\data[0][12] ) );
  DFFSR \data_reg[0][11]  ( .D(\nxt_data[0][11] ), .CLK(clk), .R(n210), .S(
        1'b1), .Q(\data[0][11] ) );
  DFFSR \data_reg[0][10]  ( .D(\nxt_data[0][10] ), .CLK(clk), .R(n210), .S(
        1'b1), .Q(\data[0][10] ) );
  DFFSR \data_reg[0][9]  ( .D(\nxt_data[0][9] ), .CLK(clk), .R(n210), .S(1'b1), 
        .Q(\data[0][9] ) );
  DFFSR \data_reg[0][8]  ( .D(\nxt_data[0][8] ), .CLK(clk), .R(n210), .S(1'b1), 
        .Q(\data[0][8] ) );
  DFFSR \data_reg[0][7]  ( .D(\nxt_data[0][7] ), .CLK(clk), .R(n210), .S(1'b1), 
        .Q(\data[0][7] ) );
  DFFSR \data_reg[0][6]  ( .D(\nxt_data[0][6] ), .CLK(clk), .R(n210), .S(1'b1), 
        .Q(\data[0][6] ) );
  DFFSR \data_reg[0][5]  ( .D(\nxt_data[0][5] ), .CLK(clk), .R(n210), .S(1'b1), 
        .Q(\data[0][5] ) );
  DFFSR \data_reg[0][4]  ( .D(\nxt_data[0][4] ), .CLK(clk), .R(n210), .S(1'b1), 
        .Q(\data[0][4] ) );
  DFFSR \data_reg[0][3]  ( .D(\nxt_data[0][3] ), .CLK(clk), .R(n210), .S(1'b1), 
        .Q(\data[0][3] ) );
  DFFSR \data_reg[0][2]  ( .D(\nxt_data[0][2] ), .CLK(clk), .R(n210), .S(1'b1), 
        .Q(\data[0][2] ) );
  DFFSR \data_reg[0][1]  ( .D(\nxt_data[0][1] ), .CLK(clk), .R(n210), .S(1'b1), 
        .Q(\data[0][1] ) );
  DFFSR \data_reg[0][0]  ( .D(\nxt_data[0][0] ), .CLK(clk), .R(n210), .S(1'b1), 
        .Q(\data[0][0] ) );
  flex_indexer_NUM_CNT_BITS2_1 Write_pointer ( .clk(clk), .n_rst(n210), 
        .clear(1'b0), .count_enable(n387), .rollover_val({1'b1, 1'b1}), 
        .count_out(w_pointer) );
  flex_indexer_NUM_CNT_BITS2_0 Read_pointer ( .clk(clk), .n_rst(n210), .clear(
        1'b0), .count_enable(_2_net_), .rollover_val({1'b1, 1'b1}), 
        .count_out({N5, N4}) );
  INVX2 U131 ( .A(n205), .Y(n203) );
  INVX8 U132 ( .A(n205), .Y(n2) );
  AND2X2 U133 ( .A(net5035), .B(net5180), .Y(n1) );
  INVX1 U134 ( .A(net5101), .Y(net5099) );
  INVX2 U135 ( .A(n209), .Y(n3) );
  INVX4 U136 ( .A(net5158), .Y(n4) );
  INVX4 U137 ( .A(net5158), .Y(n5) );
  INVX4 U138 ( .A(net5158), .Y(net5123) );
  INVX4 U139 ( .A(net5160), .Y(n6) );
  INVX4 U140 ( .A(net5160), .Y(n7) );
  INVX4 U141 ( .A(net5160), .Y(net5121) );
  XOR2X1 U142 ( .A(N4), .B(net5201), .Y(net5842) );
  BUFX4 U143 ( .A(w_pointer[0]), .Y(net5201) );
  NAND2X1 U144 ( .A(net5036), .B(net5842), .Y(net5211) );
  NOR2X1 U145 ( .A(net5201), .B(net4965), .Y(net5035) );
  XOR2X1 U146 ( .A(net5201), .B(N4), .Y(net5037) );
  AND2X2 U147 ( .A(n1), .B(net5211), .Y(n8) );
  INVX2 U148 ( .A(w_enable), .Y(net4965) );
  BUFX2 U149 ( .A(net5191), .Y(net5180) );
  INVX4 U150 ( .A(n8), .Y(net5133) );
  XOR2X1 U151 ( .A(net5841), .B(N5), .Y(net5036) );
  INVX1 U152 ( .A(net5211), .Y(net2542) );
  NAND3X1 U153 ( .A(net5000), .B(net5180), .C(net5211), .Y(net4999) );
  MUX2X1 U154 ( .B(n137), .A(net4924), .S(net5127), .Y(\nxt_data[0][0] ) );
  INVX2 U155 ( .A(\data[0][0] ), .Y(n137) );
  INVX2 U156 ( .A(w_data[0]), .Y(net4924) );
  INVX8 U157 ( .A(net5133), .Y(net5127) );
  INVX8 U158 ( .A(net5133), .Y(net5129) );
  XOR2X1 U159 ( .A(net4928), .B(w_pointer[0]), .Y(net5841) );
  INVX2 U160 ( .A(w_pointer[1]), .Y(net4928) );
  INVX1 U161 ( .A(N4), .Y(net5079) );
  BUFX2 U162 ( .A(N4), .Y(\C447/net5073 ) );
  BUFX2 U163 ( .A(N4), .Y(\C447/net5071 ) );
  BUFX2 U164 ( .A(N4), .Y(\C447/net5069 ) );
  BUFX2 U165 ( .A(N4), .Y(\C447/net5067 ) );
  BUFX2 U166 ( .A(N4), .Y(\C447/net5075 ) );
  INVX2 U167 ( .A(\C447/net5091 ), .Y(\C447/net5087 ) );
  INVX2 U168 ( .A(net5099), .Y(\C447/net5091 ) );
  XNOR2X1 U169 ( .A(net5101), .B(net5191), .Y(n217) );
  BUFX2 U170 ( .A(n_rst), .Y(n215) );
  MUX2X1 U171 ( .B(n138), .A(n139), .S(net5099), .Y(r_data[0]) );
  MUX2X1 U172 ( .B(n140), .A(n141), .S(net5099), .Y(r_data[1]) );
  MUX2X1 U173 ( .B(n142), .A(n143), .S(net5099), .Y(r_data[2]) );
  MUX2X1 U174 ( .B(n144), .A(n145), .S(net5099), .Y(r_data[3]) );
  MUX2X1 U175 ( .B(n146), .A(n147), .S(net5099), .Y(r_data[4]) );
  MUX2X1 U176 ( .B(n148), .A(n149), .S(net5099), .Y(r_data[5]) );
  MUX2X1 U177 ( .B(n150), .A(n151), .S(\C447/net5087 ), .Y(r_data[6]) );
  MUX2X1 U178 ( .B(n152), .A(n153), .S(\C447/net5087 ), .Y(r_data[7]) );
  MUX2X1 U179 ( .B(n154), .A(n155), .S(\C447/net5087 ), .Y(r_data[8]) );
  MUX2X1 U180 ( .B(n156), .A(n157), .S(\C447/net5087 ), .Y(r_data[9]) );
  MUX2X1 U181 ( .B(n158), .A(n159), .S(\C447/net5087 ), .Y(r_data[10]) );
  MUX2X1 U182 ( .B(n160), .A(n161), .S(\C447/net5087 ), .Y(r_data[11]) );
  MUX2X1 U183 ( .B(n162), .A(n163), .S(\C447/net5087 ), .Y(r_data[12]) );
  MUX2X1 U184 ( .B(n164), .A(n165), .S(\C447/net5087 ), .Y(r_data[13]) );
  MUX2X1 U185 ( .B(n166), .A(n167), .S(\C447/net5087 ), .Y(r_data[14]) );
  MUX2X1 U186 ( .B(n168), .A(n169), .S(\C447/net5087 ), .Y(r_data[15]) );
  MUX2X1 U187 ( .B(n170), .A(n171), .S(\C447/net5087 ), .Y(r_data[16]) );
  MUX2X1 U188 ( .B(n172), .A(n173), .S(\C447/net5087 ), .Y(r_data[17]) );
  MUX2X1 U189 ( .B(n174), .A(n175), .S(\C447/net5087 ), .Y(r_data[18]) );
  MUX2X1 U190 ( .B(n176), .A(n177), .S(net5099), .Y(r_data[19]) );
  MUX2X1 U191 ( .B(n178), .A(n179), .S(net5099), .Y(r_data[20]) );
  MUX2X1 U192 ( .B(n180), .A(n181), .S(net5099), .Y(r_data[21]) );
  MUX2X1 U193 ( .B(n182), .A(n183), .S(net5099), .Y(r_data[22]) );
  MUX2X1 U194 ( .B(n184), .A(n185), .S(\C447/net5087 ), .Y(r_data[23]) );
  MUX2X1 U195 ( .B(n186), .A(n187), .S(\C447/net5087 ), .Y(r_data[24]) );
  MUX2X1 U196 ( .B(n188), .A(n189), .S(\C447/net5087 ), .Y(r_data[25]) );
  MUX2X1 U197 ( .B(n190), .A(n191), .S(\C447/net5087 ), .Y(r_data[26]) );
  MUX2X1 U198 ( .B(n192), .A(n193), .S(\C447/net5087 ), .Y(r_data[27]) );
  MUX2X1 U199 ( .B(n194), .A(n195), .S(\C447/net5087 ), .Y(r_data[28]) );
  MUX2X1 U200 ( .B(n196), .A(n197), .S(\C447/net5087 ), .Y(r_data[29]) );
  MUX2X1 U201 ( .B(n198), .A(n199), .S(\C447/net5087 ), .Y(r_data[30]) );
  MUX2X1 U202 ( .B(n200), .A(n201), .S(\C447/net5087 ), .Y(r_data[31]) );
  MUX2X1 U203 ( .B(\data[2][0] ), .A(\data[3][0] ), .S(\C447/net5075 ), .Y(
        n139) );
  MUX2X1 U204 ( .B(\data[0][0] ), .A(\data[1][0] ), .S(\C447/net5075 ), .Y(
        n138) );
  MUX2X1 U205 ( .B(\data[2][1] ), .A(\data[3][1] ), .S(\C447/net5075 ), .Y(
        n141) );
  MUX2X1 U206 ( .B(\data[0][1] ), .A(\data[1][1] ), .S(\C447/net5075 ), .Y(
        n140) );
  MUX2X1 U207 ( .B(\data[2][2] ), .A(\data[3][2] ), .S(\C447/net5075 ), .Y(
        n143) );
  MUX2X1 U208 ( .B(\data[0][2] ), .A(\data[1][2] ), .S(\C447/net5075 ), .Y(
        n142) );
  MUX2X1 U209 ( .B(\data[2][3] ), .A(\data[3][3] ), .S(\C447/net5075 ), .Y(
        n145) );
  MUX2X1 U210 ( .B(\data[0][3] ), .A(\data[1][3] ), .S(\C447/net5075 ), .Y(
        n144) );
  MUX2X1 U211 ( .B(\data[2][4] ), .A(\data[3][4] ), .S(\C447/net5075 ), .Y(
        n147) );
  MUX2X1 U212 ( .B(\data[0][4] ), .A(\data[1][4] ), .S(\C447/net5075 ), .Y(
        n146) );
  MUX2X1 U213 ( .B(\data[2][5] ), .A(\data[3][5] ), .S(\C447/net5075 ), .Y(
        n149) );
  MUX2X1 U214 ( .B(\data[0][5] ), .A(\data[1][5] ), .S(\C447/net5075 ), .Y(
        n148) );
  MUX2X1 U215 ( .B(\data[2][6] ), .A(\data[3][6] ), .S(\C447/net5073 ), .Y(
        n151) );
  MUX2X1 U216 ( .B(\data[0][6] ), .A(\data[1][6] ), .S(\C447/net5073 ), .Y(
        n150) );
  MUX2X1 U217 ( .B(\data[2][7] ), .A(\data[3][7] ), .S(\C447/net5073 ), .Y(
        n153) );
  MUX2X1 U218 ( .B(\data[0][7] ), .A(\data[1][7] ), .S(\C447/net5073 ), .Y(
        n152) );
  MUX2X1 U219 ( .B(\data[2][8] ), .A(\data[3][8] ), .S(\C447/net5073 ), .Y(
        n155) );
  MUX2X1 U220 ( .B(\data[0][8] ), .A(\data[1][8] ), .S(\C447/net5073 ), .Y(
        n154) );
  MUX2X1 U221 ( .B(\data[2][9] ), .A(\data[3][9] ), .S(\C447/net5073 ), .Y(
        n157) );
  MUX2X1 U222 ( .B(\data[0][9] ), .A(\data[1][9] ), .S(\C447/net5073 ), .Y(
        n156) );
  MUX2X1 U223 ( .B(\data[2][10] ), .A(\data[3][10] ), .S(\C447/net5073 ), .Y(
        n159) );
  MUX2X1 U224 ( .B(\data[0][10] ), .A(\data[1][10] ), .S(\C447/net5073 ), .Y(
        n158) );
  MUX2X1 U225 ( .B(\data[2][11] ), .A(\data[3][11] ), .S(\C447/net5073 ), .Y(
        n161) );
  MUX2X1 U226 ( .B(\data[0][11] ), .A(\data[1][11] ), .S(\C447/net5073 ), .Y(
        n160) );
  MUX2X1 U227 ( .B(\data[2][12] ), .A(\data[3][12] ), .S(\C447/net5073 ), .Y(
        n163) );
  MUX2X1 U228 ( .B(\data[0][12] ), .A(\data[1][12] ), .S(\C447/net5071 ), .Y(
        n162) );
  MUX2X1 U229 ( .B(\data[2][13] ), .A(\data[3][13] ), .S(\C447/net5071 ), .Y(
        n165) );
  MUX2X1 U230 ( .B(\data[0][13] ), .A(\data[1][13] ), .S(\C447/net5071 ), .Y(
        n164) );
  MUX2X1 U231 ( .B(\data[2][14] ), .A(\data[3][14] ), .S(\C447/net5071 ), .Y(
        n167) );
  MUX2X1 U232 ( .B(\data[0][14] ), .A(\data[1][14] ), .S(\C447/net5071 ), .Y(
        n166) );
  MUX2X1 U233 ( .B(\data[2][15] ), .A(\data[3][15] ), .S(\C447/net5071 ), .Y(
        n169) );
  MUX2X1 U234 ( .B(\data[0][15] ), .A(\data[1][15] ), .S(\C447/net5071 ), .Y(
        n168) );
  MUX2X1 U235 ( .B(\data[2][16] ), .A(\data[3][16] ), .S(\C447/net5071 ), .Y(
        n171) );
  MUX2X1 U236 ( .B(\data[0][16] ), .A(\data[1][16] ), .S(\C447/net5071 ), .Y(
        n170) );
  MUX2X1 U237 ( .B(\data[2][17] ), .A(\data[3][17] ), .S(\C447/net5071 ), .Y(
        n173) );
  MUX2X1 U238 ( .B(\data[0][17] ), .A(\data[1][17] ), .S(\C447/net5071 ), .Y(
        n172) );
  MUX2X1 U239 ( .B(\data[2][18] ), .A(\data[3][18] ), .S(\C447/net5071 ), .Y(
        n175) );
  MUX2X1 U240 ( .B(\data[0][18] ), .A(\data[1][18] ), .S(\C447/net5071 ), .Y(
        n174) );
  MUX2X1 U241 ( .B(\data[2][19] ), .A(\data[3][19] ), .S(\C447/net5069 ), .Y(
        n177) );
  MUX2X1 U242 ( .B(\data[0][19] ), .A(\data[1][19] ), .S(\C447/net5069 ), .Y(
        n176) );
  MUX2X1 U243 ( .B(\data[2][20] ), .A(\data[3][20] ), .S(\C447/net5069 ), .Y(
        n179) );
  MUX2X1 U244 ( .B(\data[0][20] ), .A(\data[1][20] ), .S(\C447/net5069 ), .Y(
        n178) );
  MUX2X1 U245 ( .B(\data[2][21] ), .A(\data[3][21] ), .S(\C447/net5069 ), .Y(
        n181) );
  MUX2X1 U246 ( .B(\data[0][21] ), .A(\data[1][21] ), .S(\C447/net5069 ), .Y(
        n180) );
  MUX2X1 U247 ( .B(\data[2][22] ), .A(\data[3][22] ), .S(\C447/net5069 ), .Y(
        n183) );
  MUX2X1 U248 ( .B(\data[0][22] ), .A(\data[1][22] ), .S(\C447/net5069 ), .Y(
        n182) );
  MUX2X1 U249 ( .B(\data[2][23] ), .A(\data[3][23] ), .S(\C447/net5069 ), .Y(
        n185) );
  MUX2X1 U250 ( .B(\data[0][23] ), .A(\data[1][23] ), .S(\C447/net5069 ), .Y(
        n184) );
  MUX2X1 U251 ( .B(\data[2][24] ), .A(\data[3][24] ), .S(\C447/net5069 ), .Y(
        n187) );
  MUX2X1 U252 ( .B(\data[0][24] ), .A(\data[1][24] ), .S(\C447/net5069 ), .Y(
        n186) );
  MUX2X1 U253 ( .B(\data[2][25] ), .A(\data[3][25] ), .S(\C447/net5069 ), .Y(
        n189) );
  MUX2X1 U254 ( .B(\data[0][25] ), .A(\data[1][25] ), .S(\C447/net5067 ), .Y(
        n188) );
  MUX2X1 U255 ( .B(\data[2][26] ), .A(\data[3][26] ), .S(\C447/net5067 ), .Y(
        n191) );
  MUX2X1 U256 ( .B(\data[0][26] ), .A(\data[1][26] ), .S(\C447/net5067 ), .Y(
        n190) );
  MUX2X1 U257 ( .B(\data[2][27] ), .A(\data[3][27] ), .S(\C447/net5067 ), .Y(
        n193) );
  MUX2X1 U258 ( .B(\data[0][27] ), .A(\data[1][27] ), .S(\C447/net5067 ), .Y(
        n192) );
  MUX2X1 U259 ( .B(\data[2][28] ), .A(\data[3][28] ), .S(\C447/net5067 ), .Y(
        n195) );
  MUX2X1 U260 ( .B(\data[0][28] ), .A(\data[1][28] ), .S(\C447/net5067 ), .Y(
        n194) );
  MUX2X1 U261 ( .B(\data[2][29] ), .A(\data[3][29] ), .S(\C447/net5067 ), .Y(
        n197) );
  MUX2X1 U262 ( .B(\data[0][29] ), .A(\data[1][29] ), .S(\C447/net5067 ), .Y(
        n196) );
  MUX2X1 U263 ( .B(\data[2][30] ), .A(\data[3][30] ), .S(\C447/net5067 ), .Y(
        n199) );
  MUX2X1 U264 ( .B(\data[0][30] ), .A(\data[1][30] ), .S(\C447/net5067 ), .Y(
        n198) );
  MUX2X1 U265 ( .B(\data[2][31] ), .A(\data[3][31] ), .S(\C447/net5067 ), .Y(
        n201) );
  MUX2X1 U266 ( .B(\data[0][31] ), .A(\data[1][31] ), .S(\C447/net5067 ), .Y(
        n200) );
  INVX4 U267 ( .A(n322), .Y(n384) );
  INVX8 U268 ( .A(n384), .Y(n209) );
  INVX4 U269 ( .A(N5), .Y(net5101) );
  INVX1 U270 ( .A(net4929), .Y(net5196) );
  INVX1 U271 ( .A(w_pointer[1]), .Y(net5191) );
  INVX1 U272 ( .A(net4928), .Y(net5185) );
  INVX1 U273 ( .A(net5185), .Y(net5186) );
  BUFX4 U274 ( .A(net4999), .Y(net5160) );
  BUFX4 U275 ( .A(net4999), .Y(net5158) );
  INVX4 U276 ( .A(n205), .Y(n204) );
  INVX4 U277 ( .A(n286), .Y(n318) );
  INVX4 U278 ( .A(n209), .Y(n208) );
  INVX8 U279 ( .A(n205), .Y(n202) );
  INVX8 U280 ( .A(n318), .Y(n205) );
  INVX8 U281 ( .A(n209), .Y(n206) );
  INVX8 U282 ( .A(n209), .Y(n207) );
  BUFX4 U283 ( .A(n_rst), .Y(n210) );
  BUFX4 U284 ( .A(n_rst), .Y(n211) );
  BUFX4 U285 ( .A(n_rst), .Y(n212) );
  BUFX4 U286 ( .A(n_rst), .Y(n213) );
  BUFX4 U287 ( .A(n_rst), .Y(n214) );
  INVX2 U288 ( .A(w_pointer[0]), .Y(net4929) );
  XOR2X1 U289 ( .A(net4929), .B(N4), .Y(n216) );
  NAND2X1 U290 ( .A(n216), .B(n217), .Y(n221) );
  AND2X2 U291 ( .A(r_enable), .B(n221), .Y(_2_net_) );
  NOR2X1 U292 ( .A(net4929), .B(n217), .Y(n220) );
  NAND2X1 U293 ( .A(N4), .B(n217), .Y(n218) );
  OAI21X1 U294 ( .A(net5196), .B(n218), .C(w_enable), .Y(n219) );
  AOI21X1 U295 ( .A(n220), .B(net5079), .C(n219), .Y(n387) );
  INVX2 U296 ( .A(n221), .Y(N14) );
  NAND2X1 U297 ( .A(net5036), .B(net5037), .Y(n320) );
  INVX2 U298 ( .A(\data[0][1] ), .Y(n222) );
  INVX2 U299 ( .A(w_data[1]), .Y(n324) );
  MUX2X1 U300 ( .B(n222), .A(n324), .S(net5127), .Y(\nxt_data[0][1] ) );
  INVX2 U301 ( .A(\data[0][2] ), .Y(n223) );
  INVX2 U302 ( .A(w_data[2]), .Y(n326) );
  MUX2X1 U303 ( .B(n223), .A(n326), .S(net5127), .Y(\nxt_data[0][2] ) );
  INVX2 U304 ( .A(\data[0][3] ), .Y(n224) );
  INVX2 U305 ( .A(w_data[3]), .Y(n328) );
  MUX2X1 U306 ( .B(n224), .A(n328), .S(net5127), .Y(\nxt_data[0][3] ) );
  INVX2 U307 ( .A(\data[0][4] ), .Y(n225) );
  INVX2 U308 ( .A(w_data[4]), .Y(n330) );
  MUX2X1 U309 ( .B(n225), .A(n330), .S(net5127), .Y(\nxt_data[0][4] ) );
  INVX2 U310 ( .A(\data[0][5] ), .Y(n226) );
  INVX2 U311 ( .A(w_data[5]), .Y(n332) );
  MUX2X1 U312 ( .B(n226), .A(n332), .S(net5127), .Y(\nxt_data[0][5] ) );
  INVX2 U313 ( .A(\data[0][6] ), .Y(n227) );
  INVX2 U314 ( .A(w_data[6]), .Y(n334) );
  MUX2X1 U315 ( .B(n227), .A(n334), .S(net5127), .Y(\nxt_data[0][6] ) );
  INVX2 U316 ( .A(\data[0][7] ), .Y(n228) );
  INVX2 U317 ( .A(w_data[7]), .Y(n336) );
  MUX2X1 U318 ( .B(n228), .A(n336), .S(net5127), .Y(\nxt_data[0][7] ) );
  INVX2 U319 ( .A(\data[0][8] ), .Y(n229) );
  INVX2 U320 ( .A(w_data[8]), .Y(n338) );
  MUX2X1 U321 ( .B(n229), .A(n338), .S(net5127), .Y(\nxt_data[0][8] ) );
  INVX2 U322 ( .A(\data[0][9] ), .Y(n230) );
  INVX2 U323 ( .A(w_data[9]), .Y(n340) );
  MUX2X1 U324 ( .B(n230), .A(n340), .S(net5127), .Y(\nxt_data[0][9] ) );
  INVX2 U325 ( .A(\data[0][10] ), .Y(n231) );
  INVX2 U326 ( .A(w_data[10]), .Y(n342) );
  MUX2X1 U327 ( .B(n231), .A(n342), .S(net5127), .Y(\nxt_data[0][10] ) );
  INVX2 U328 ( .A(\data[0][11] ), .Y(n232) );
  INVX2 U329 ( .A(w_data[11]), .Y(n344) );
  MUX2X1 U330 ( .B(n232), .A(n344), .S(net5127), .Y(\nxt_data[0][11] ) );
  INVX2 U331 ( .A(\data[0][12] ), .Y(n233) );
  INVX2 U332 ( .A(w_data[12]), .Y(n346) );
  MUX2X1 U333 ( .B(n233), .A(n346), .S(net5127), .Y(\nxt_data[0][12] ) );
  INVX2 U334 ( .A(\data[0][13] ), .Y(n234) );
  INVX2 U335 ( .A(w_data[13]), .Y(n348) );
  MUX2X1 U336 ( .B(n234), .A(n348), .S(net5129), .Y(\nxt_data[0][13] ) );
  INVX2 U337 ( .A(\data[0][14] ), .Y(n235) );
  INVX2 U338 ( .A(w_data[14]), .Y(n350) );
  MUX2X1 U339 ( .B(n235), .A(n350), .S(net5129), .Y(\nxt_data[0][14] ) );
  INVX2 U340 ( .A(\data[0][15] ), .Y(n236) );
  INVX2 U341 ( .A(w_data[15]), .Y(n352) );
  MUX2X1 U342 ( .B(n236), .A(n352), .S(net5129), .Y(\nxt_data[0][15] ) );
  INVX2 U343 ( .A(\data[0][16] ), .Y(n237) );
  INVX2 U344 ( .A(w_data[16]), .Y(n354) );
  MUX2X1 U345 ( .B(n237), .A(n354), .S(net5129), .Y(\nxt_data[0][16] ) );
  INVX2 U346 ( .A(\data[0][17] ), .Y(n238) );
  INVX2 U347 ( .A(w_data[17]), .Y(n356) );
  MUX2X1 U348 ( .B(n238), .A(n356), .S(net5129), .Y(\nxt_data[0][17] ) );
  INVX2 U349 ( .A(\data[0][18] ), .Y(n239) );
  INVX2 U350 ( .A(w_data[18]), .Y(n358) );
  MUX2X1 U351 ( .B(n239), .A(n358), .S(net5129), .Y(\nxt_data[0][18] ) );
  INVX2 U352 ( .A(\data[0][19] ), .Y(n240) );
  INVX2 U353 ( .A(w_data[19]), .Y(n360) );
  MUX2X1 U354 ( .B(n240), .A(n360), .S(net5129), .Y(\nxt_data[0][19] ) );
  INVX2 U355 ( .A(\data[0][20] ), .Y(n241) );
  INVX2 U356 ( .A(w_data[20]), .Y(n362) );
  MUX2X1 U357 ( .B(n241), .A(n362), .S(net5129), .Y(\nxt_data[0][20] ) );
  INVX2 U358 ( .A(\data[0][21] ), .Y(n242) );
  INVX2 U359 ( .A(w_data[21]), .Y(n364) );
  MUX2X1 U360 ( .B(n242), .A(n364), .S(net5129), .Y(\nxt_data[0][21] ) );
  INVX2 U361 ( .A(\data[0][22] ), .Y(n243) );
  INVX2 U362 ( .A(w_data[22]), .Y(n366) );
  MUX2X1 U363 ( .B(n243), .A(n366), .S(net5129), .Y(\nxt_data[0][22] ) );
  INVX2 U364 ( .A(\data[0][23] ), .Y(n244) );
  INVX2 U365 ( .A(w_data[23]), .Y(n368) );
  MUX2X1 U366 ( .B(n244), .A(n368), .S(net5129), .Y(\nxt_data[0][23] ) );
  INVX2 U367 ( .A(\data[0][24] ), .Y(n245) );
  INVX2 U368 ( .A(w_data[24]), .Y(n370) );
  MUX2X1 U369 ( .B(n245), .A(n370), .S(net5129), .Y(\nxt_data[0][24] ) );
  INVX2 U370 ( .A(\data[0][25] ), .Y(n246) );
  INVX2 U371 ( .A(w_data[25]), .Y(n372) );
  MUX2X1 U372 ( .B(n246), .A(n372), .S(net5129), .Y(\nxt_data[0][25] ) );
  INVX2 U373 ( .A(\data[0][26] ), .Y(n247) );
  INVX2 U374 ( .A(w_data[26]), .Y(n374) );
  MUX2X1 U375 ( .B(n247), .A(n374), .S(net5127), .Y(\nxt_data[0][26] ) );
  INVX2 U376 ( .A(\data[0][27] ), .Y(n248) );
  INVX2 U377 ( .A(w_data[27]), .Y(n376) );
  MUX2X1 U378 ( .B(n248), .A(n376), .S(net5129), .Y(\nxt_data[0][27] ) );
  INVX2 U379 ( .A(\data[0][28] ), .Y(n249) );
  INVX2 U380 ( .A(w_data[28]), .Y(n378) );
  MUX2X1 U381 ( .B(n249), .A(n378), .S(net5127), .Y(\nxt_data[0][28] ) );
  INVX2 U382 ( .A(\data[0][29] ), .Y(n250) );
  INVX2 U383 ( .A(w_data[29]), .Y(n380) );
  MUX2X1 U384 ( .B(n250), .A(n380), .S(net5127), .Y(\nxt_data[0][29] ) );
  INVX2 U385 ( .A(\data[0][30] ), .Y(n251) );
  INVX2 U386 ( .A(w_data[30]), .Y(n382) );
  MUX2X1 U387 ( .B(n251), .A(n382), .S(net5129), .Y(\nxt_data[0][30] ) );
  INVX2 U388 ( .A(\data[0][31] ), .Y(n252) );
  INVX2 U389 ( .A(w_data[31]), .Y(n385) );
  MUX2X1 U390 ( .B(n252), .A(n385), .S(net5129), .Y(\nxt_data[0][31] ) );
  INVX2 U391 ( .A(\data[1][0] ), .Y(n253) );
  NOR2X1 U392 ( .A(net4929), .B(net4965), .Y(net5000) );
  MUX2X1 U393 ( .B(n253), .A(net4924), .S(net5121), .Y(\nxt_data[1][0] ) );
  INVX2 U394 ( .A(\data[1][1] ), .Y(n254) );
  MUX2X1 U395 ( .B(n254), .A(n324), .S(net5123), .Y(\nxt_data[1][1] ) );
  INVX2 U396 ( .A(\data[1][2] ), .Y(n255) );
  MUX2X1 U397 ( .B(n255), .A(n326), .S(net5121), .Y(\nxt_data[1][2] ) );
  INVX2 U398 ( .A(\data[1][3] ), .Y(n256) );
  MUX2X1 U399 ( .B(n256), .A(n328), .S(net5123), .Y(\nxt_data[1][3] ) );
  INVX2 U400 ( .A(\data[1][4] ), .Y(n257) );
  MUX2X1 U401 ( .B(n257), .A(n330), .S(net5123), .Y(\nxt_data[1][4] ) );
  INVX2 U402 ( .A(\data[1][5] ), .Y(n258) );
  MUX2X1 U403 ( .B(n258), .A(n332), .S(net5123), .Y(\nxt_data[1][5] ) );
  INVX2 U404 ( .A(\data[1][6] ), .Y(n259) );
  MUX2X1 U405 ( .B(n259), .A(n334), .S(net5123), .Y(\nxt_data[1][6] ) );
  INVX2 U406 ( .A(\data[1][7] ), .Y(n260) );
  MUX2X1 U407 ( .B(n260), .A(n336), .S(n5), .Y(\nxt_data[1][7] ) );
  INVX2 U408 ( .A(\data[1][8] ), .Y(n261) );
  MUX2X1 U409 ( .B(n261), .A(n338), .S(net5121), .Y(\nxt_data[1][8] ) );
  INVX2 U410 ( .A(\data[1][9] ), .Y(n262) );
  MUX2X1 U411 ( .B(n262), .A(n340), .S(net5123), .Y(\nxt_data[1][9] ) );
  INVX2 U412 ( .A(\data[1][10] ), .Y(n263) );
  MUX2X1 U413 ( .B(n263), .A(n342), .S(n4), .Y(\nxt_data[1][10] ) );
  INVX2 U414 ( .A(\data[1][11] ), .Y(n264) );
  MUX2X1 U415 ( .B(n264), .A(n344), .S(n5), .Y(\nxt_data[1][11] ) );
  INVX2 U416 ( .A(\data[1][12] ), .Y(n265) );
  MUX2X1 U417 ( .B(n265), .A(n346), .S(n4), .Y(\nxt_data[1][12] ) );
  INVX2 U418 ( .A(\data[1][13] ), .Y(n266) );
  MUX2X1 U419 ( .B(n266), .A(n348), .S(n6), .Y(\nxt_data[1][13] ) );
  INVX2 U420 ( .A(\data[1][14] ), .Y(n267) );
  MUX2X1 U421 ( .B(n267), .A(n350), .S(n7), .Y(\nxt_data[1][14] ) );
  INVX2 U422 ( .A(\data[1][15] ), .Y(n268) );
  MUX2X1 U423 ( .B(n268), .A(n352), .S(n6), .Y(\nxt_data[1][15] ) );
  INVX2 U424 ( .A(\data[1][16] ), .Y(n269) );
  MUX2X1 U425 ( .B(n269), .A(n354), .S(n7), .Y(\nxt_data[1][16] ) );
  INVX2 U426 ( .A(\data[1][17] ), .Y(n270) );
  MUX2X1 U427 ( .B(n270), .A(n356), .S(n6), .Y(\nxt_data[1][17] ) );
  INVX2 U428 ( .A(\data[1][18] ), .Y(n271) );
  MUX2X1 U429 ( .B(n271), .A(n358), .S(n7), .Y(\nxt_data[1][18] ) );
  INVX2 U430 ( .A(\data[1][19] ), .Y(n272) );
  MUX2X1 U431 ( .B(n272), .A(n360), .S(n6), .Y(\nxt_data[1][19] ) );
  INVX2 U432 ( .A(\data[1][20] ), .Y(n273) );
  MUX2X1 U433 ( .B(n273), .A(n362), .S(n7), .Y(\nxt_data[1][20] ) );
  INVX2 U434 ( .A(\data[1][21] ), .Y(n274) );
  MUX2X1 U435 ( .B(n274), .A(n364), .S(n6), .Y(\nxt_data[1][21] ) );
  INVX2 U436 ( .A(\data[1][22] ), .Y(n275) );
  MUX2X1 U437 ( .B(n275), .A(n366), .S(n7), .Y(\nxt_data[1][22] ) );
  INVX2 U438 ( .A(\data[1][23] ), .Y(n276) );
  MUX2X1 U439 ( .B(n276), .A(n368), .S(net5121), .Y(\nxt_data[1][23] ) );
  INVX2 U440 ( .A(\data[1][24] ), .Y(n277) );
  MUX2X1 U441 ( .B(n277), .A(n370), .S(net5121), .Y(\nxt_data[1][24] ) );
  INVX2 U442 ( .A(\data[1][25] ), .Y(n278) );
  MUX2X1 U443 ( .B(n278), .A(n372), .S(net5121), .Y(\nxt_data[1][25] ) );
  INVX2 U444 ( .A(\data[1][26] ), .Y(n279) );
  MUX2X1 U445 ( .B(n279), .A(n374), .S(n4), .Y(\nxt_data[1][26] ) );
  INVX2 U446 ( .A(\data[1][27] ), .Y(n280) );
  MUX2X1 U447 ( .B(n280), .A(n376), .S(n5), .Y(\nxt_data[1][27] ) );
  INVX2 U448 ( .A(\data[1][28] ), .Y(n281) );
  MUX2X1 U449 ( .B(n281), .A(n378), .S(n4), .Y(\nxt_data[1][28] ) );
  INVX2 U450 ( .A(\data[1][29] ), .Y(n282) );
  MUX2X1 U451 ( .B(n282), .A(n380), .S(n5), .Y(\nxt_data[1][29] ) );
  INVX2 U452 ( .A(\data[1][30] ), .Y(n283) );
  MUX2X1 U453 ( .B(n283), .A(n382), .S(n4), .Y(\nxt_data[1][30] ) );
  INVX2 U454 ( .A(\data[1][31] ), .Y(n284) );
  MUX2X1 U455 ( .B(n284), .A(n385), .S(n5), .Y(\nxt_data[1][31] ) );
  INVX2 U456 ( .A(\data[2][0] ), .Y(n287) );
  NOR2X1 U457 ( .A(net5186), .B(net4965), .Y(n285) );
  NAND3X1 U458 ( .A(n285), .B(net4929), .C(n320), .Y(n286) );
  MUX2X1 U459 ( .B(n287), .A(net4924), .S(n202), .Y(\nxt_data[2][0] ) );
  INVX2 U460 ( .A(\data[2][1] ), .Y(n288) );
  MUX2X1 U461 ( .B(n288), .A(n324), .S(n202), .Y(\nxt_data[2][1] ) );
  INVX2 U462 ( .A(\data[2][2] ), .Y(n289) );
  MUX2X1 U463 ( .B(n289), .A(n326), .S(n202), .Y(\nxt_data[2][2] ) );
  INVX2 U464 ( .A(\data[2][3] ), .Y(n290) );
  MUX2X1 U465 ( .B(n290), .A(n328), .S(n202), .Y(\nxt_data[2][3] ) );
  INVX2 U466 ( .A(\data[2][4] ), .Y(n291) );
  MUX2X1 U467 ( .B(n291), .A(n330), .S(n202), .Y(\nxt_data[2][4] ) );
  INVX2 U468 ( .A(\data[2][5] ), .Y(n292) );
  MUX2X1 U469 ( .B(n292), .A(n332), .S(n202), .Y(\nxt_data[2][5] ) );
  INVX2 U470 ( .A(\data[2][6] ), .Y(n293) );
  MUX2X1 U471 ( .B(n293), .A(n334), .S(n202), .Y(\nxt_data[2][6] ) );
  INVX2 U472 ( .A(\data[2][7] ), .Y(n294) );
  MUX2X1 U473 ( .B(n294), .A(n336), .S(n202), .Y(\nxt_data[2][7] ) );
  INVX2 U474 ( .A(\data[2][8] ), .Y(n295) );
  MUX2X1 U475 ( .B(n295), .A(n338), .S(n202), .Y(\nxt_data[2][8] ) );
  INVX2 U476 ( .A(\data[2][9] ), .Y(n296) );
  MUX2X1 U477 ( .B(n296), .A(n340), .S(n202), .Y(\nxt_data[2][9] ) );
  INVX2 U478 ( .A(\data[2][10] ), .Y(n297) );
  MUX2X1 U479 ( .B(n297), .A(n342), .S(n202), .Y(\nxt_data[2][10] ) );
  INVX2 U480 ( .A(\data[2][11] ), .Y(n298) );
  MUX2X1 U481 ( .B(n298), .A(n344), .S(n202), .Y(\nxt_data[2][11] ) );
  INVX2 U482 ( .A(\data[2][12] ), .Y(n299) );
  MUX2X1 U483 ( .B(n299), .A(n346), .S(n2), .Y(\nxt_data[2][12] ) );
  INVX2 U484 ( .A(\data[2][13] ), .Y(n300) );
  MUX2X1 U485 ( .B(n300), .A(n348), .S(n203), .Y(\nxt_data[2][13] ) );
  INVX2 U486 ( .A(\data[2][14] ), .Y(n301) );
  MUX2X1 U487 ( .B(n301), .A(n350), .S(n203), .Y(\nxt_data[2][14] ) );
  INVX2 U488 ( .A(\data[2][15] ), .Y(n302) );
  MUX2X1 U489 ( .B(n302), .A(n352), .S(n203), .Y(\nxt_data[2][15] ) );
  INVX2 U490 ( .A(\data[2][16] ), .Y(n303) );
  MUX2X1 U491 ( .B(n303), .A(n354), .S(n2), .Y(\nxt_data[2][16] ) );
  INVX2 U492 ( .A(\data[2][17] ), .Y(n304) );
  MUX2X1 U493 ( .B(n304), .A(n356), .S(n2), .Y(\nxt_data[2][17] ) );
  INVX2 U494 ( .A(\data[2][18] ), .Y(n305) );
  MUX2X1 U495 ( .B(n305), .A(n358), .S(n2), .Y(\nxt_data[2][18] ) );
  INVX2 U496 ( .A(\data[2][19] ), .Y(n306) );
  MUX2X1 U497 ( .B(n306), .A(n360), .S(n2), .Y(\nxt_data[2][19] ) );
  INVX2 U498 ( .A(\data[2][20] ), .Y(n307) );
  MUX2X1 U499 ( .B(n307), .A(n362), .S(n2), .Y(\nxt_data[2][20] ) );
  INVX2 U500 ( .A(\data[2][21] ), .Y(n308) );
  MUX2X1 U501 ( .B(n308), .A(n364), .S(n2), .Y(\nxt_data[2][21] ) );
  INVX2 U502 ( .A(\data[2][22] ), .Y(n309) );
  MUX2X1 U503 ( .B(n309), .A(n366), .S(n2), .Y(\nxt_data[2][22] ) );
  INVX2 U504 ( .A(\data[2][23] ), .Y(n310) );
  MUX2X1 U505 ( .B(n310), .A(n368), .S(n2), .Y(\nxt_data[2][23] ) );
  INVX2 U506 ( .A(\data[2][24] ), .Y(n311) );
  MUX2X1 U507 ( .B(n311), .A(n370), .S(n2), .Y(\nxt_data[2][24] ) );
  INVX2 U508 ( .A(\data[2][25] ), .Y(n312) );
  MUX2X1 U509 ( .B(n312), .A(n372), .S(n2), .Y(\nxt_data[2][25] ) );
  INVX2 U510 ( .A(\data[2][26] ), .Y(n313) );
  MUX2X1 U511 ( .B(n313), .A(n374), .S(n204), .Y(\nxt_data[2][26] ) );
  INVX2 U512 ( .A(\data[2][27] ), .Y(n314) );
  MUX2X1 U513 ( .B(n314), .A(n376), .S(n204), .Y(\nxt_data[2][27] ) );
  INVX2 U514 ( .A(\data[2][28] ), .Y(n315) );
  MUX2X1 U515 ( .B(n315), .A(n378), .S(n204), .Y(\nxt_data[2][28] ) );
  INVX2 U516 ( .A(\data[2][29] ), .Y(n316) );
  MUX2X1 U517 ( .B(n316), .A(n380), .S(n204), .Y(\nxt_data[2][29] ) );
  INVX2 U518 ( .A(\data[2][30] ), .Y(n317) );
  MUX2X1 U519 ( .B(n317), .A(n382), .S(n204), .Y(\nxt_data[2][30] ) );
  INVX2 U520 ( .A(\data[2][31] ), .Y(n319) );
  MUX2X1 U521 ( .B(n319), .A(n385), .S(n204), .Y(\nxt_data[2][31] ) );
  INVX2 U522 ( .A(\data[3][0] ), .Y(n323) );
  NOR2X1 U523 ( .A(net5180), .B(net4929), .Y(n321) );
  NAND3X1 U524 ( .A(w_enable), .B(n321), .C(n320), .Y(n322) );
  MUX2X1 U525 ( .B(n323), .A(net4924), .S(n206), .Y(\nxt_data[3][0] ) );
  INVX2 U526 ( .A(\data[3][1] ), .Y(n325) );
  MUX2X1 U527 ( .B(n325), .A(n324), .S(n206), .Y(\nxt_data[3][1] ) );
  INVX2 U528 ( .A(\data[3][2] ), .Y(n327) );
  MUX2X1 U529 ( .B(n327), .A(n326), .S(n3), .Y(\nxt_data[3][2] ) );
  INVX2 U530 ( .A(\data[3][3] ), .Y(n329) );
  MUX2X1 U531 ( .B(n329), .A(n328), .S(n206), .Y(\nxt_data[3][3] ) );
  INVX2 U532 ( .A(\data[3][4] ), .Y(n331) );
  MUX2X1 U533 ( .B(n331), .A(n330), .S(n208), .Y(\nxt_data[3][4] ) );
  INVX2 U534 ( .A(\data[3][5] ), .Y(n333) );
  MUX2X1 U535 ( .B(n333), .A(n332), .S(n206), .Y(\nxt_data[3][5] ) );
  INVX2 U536 ( .A(\data[3][6] ), .Y(n335) );
  MUX2X1 U537 ( .B(n335), .A(n334), .S(n206), .Y(\nxt_data[3][6] ) );
  INVX2 U538 ( .A(\data[3][7] ), .Y(n337) );
  MUX2X1 U539 ( .B(n337), .A(n336), .S(n3), .Y(\nxt_data[3][7] ) );
  INVX2 U540 ( .A(\data[3][8] ), .Y(n339) );
  MUX2X1 U541 ( .B(n339), .A(n338), .S(n208), .Y(\nxt_data[3][8] ) );
  INVX2 U542 ( .A(\data[3][9] ), .Y(n341) );
  MUX2X1 U543 ( .B(n341), .A(n340), .S(n206), .Y(\nxt_data[3][9] ) );
  INVX2 U544 ( .A(\data[3][10] ), .Y(n343) );
  MUX2X1 U545 ( .B(n343), .A(n342), .S(n206), .Y(\nxt_data[3][10] ) );
  INVX2 U546 ( .A(\data[3][11] ), .Y(n345) );
  MUX2X1 U547 ( .B(n345), .A(n344), .S(n208), .Y(\nxt_data[3][11] ) );
  INVX2 U548 ( .A(\data[3][12] ), .Y(n347) );
  MUX2X1 U549 ( .B(n347), .A(n346), .S(n206), .Y(\nxt_data[3][12] ) );
  INVX2 U550 ( .A(\data[3][13] ), .Y(n349) );
  MUX2X1 U551 ( .B(n349), .A(n348), .S(n208), .Y(\nxt_data[3][13] ) );
  INVX2 U552 ( .A(\data[3][14] ), .Y(n351) );
  MUX2X1 U553 ( .B(n351), .A(n350), .S(n207), .Y(\nxt_data[3][14] ) );
  INVX2 U554 ( .A(\data[3][15] ), .Y(n353) );
  MUX2X1 U555 ( .B(n353), .A(n352), .S(n207), .Y(\nxt_data[3][15] ) );
  INVX2 U556 ( .A(\data[3][16] ), .Y(n355) );
  MUX2X1 U557 ( .B(n355), .A(n354), .S(n207), .Y(\nxt_data[3][16] ) );
  INVX2 U558 ( .A(\data[3][17] ), .Y(n357) );
  MUX2X1 U559 ( .B(n357), .A(n356), .S(n207), .Y(\nxt_data[3][17] ) );
  INVX2 U560 ( .A(\data[3][18] ), .Y(n359) );
  MUX2X1 U561 ( .B(n359), .A(n358), .S(n207), .Y(\nxt_data[3][18] ) );
  INVX2 U562 ( .A(\data[3][19] ), .Y(n361) );
  MUX2X1 U563 ( .B(n361), .A(n360), .S(n207), .Y(\nxt_data[3][19] ) );
  INVX2 U564 ( .A(\data[3][20] ), .Y(n363) );
  MUX2X1 U565 ( .B(n363), .A(n362), .S(n207), .Y(\nxt_data[3][20] ) );
  INVX2 U566 ( .A(\data[3][21] ), .Y(n365) );
  MUX2X1 U567 ( .B(n365), .A(n364), .S(n207), .Y(\nxt_data[3][21] ) );
  INVX2 U568 ( .A(\data[3][22] ), .Y(n367) );
  MUX2X1 U569 ( .B(n367), .A(n366), .S(n207), .Y(\nxt_data[3][22] ) );
  INVX2 U570 ( .A(\data[3][23] ), .Y(n369) );
  MUX2X1 U571 ( .B(n369), .A(n368), .S(n207), .Y(\nxt_data[3][23] ) );
  INVX2 U572 ( .A(\data[3][24] ), .Y(n371) );
  MUX2X1 U573 ( .B(n371), .A(n370), .S(n207), .Y(\nxt_data[3][24] ) );
  INVX2 U574 ( .A(\data[3][25] ), .Y(n373) );
  MUX2X1 U575 ( .B(n373), .A(n372), .S(n207), .Y(\nxt_data[3][25] ) );
  INVX2 U576 ( .A(\data[3][26] ), .Y(n375) );
  MUX2X1 U577 ( .B(n375), .A(n374), .S(n206), .Y(\nxt_data[3][26] ) );
  INVX2 U578 ( .A(\data[3][27] ), .Y(n377) );
  MUX2X1 U579 ( .B(n377), .A(n376), .S(n3), .Y(\nxt_data[3][27] ) );
  INVX2 U580 ( .A(\data[3][28] ), .Y(n379) );
  MUX2X1 U581 ( .B(n379), .A(n378), .S(n208), .Y(\nxt_data[3][28] ) );
  INVX2 U582 ( .A(\data[3][29] ), .Y(n381) );
  MUX2X1 U583 ( .B(n381), .A(n380), .S(n206), .Y(\nxt_data[3][29] ) );
  INVX2 U584 ( .A(\data[3][30] ), .Y(n383) );
  MUX2X1 U585 ( .B(n383), .A(n382), .S(n206), .Y(\nxt_data[3][30] ) );
  INVX2 U586 ( .A(\data[3][31] ), .Y(n386) );
  MUX2X1 U587 ( .B(n386), .A(n385), .S(n208), .Y(\nxt_data[3][31] ) );
endmodule


module instruction_parser ( clk, n_rst, address_bus, data_bus, 
        read_instruction, valid_data, dependency_remove, read_data_buff, 
        read_data_enable, instruction_buffer_full, instruction_out, 
        add_instruction, out_reg, read_error, write_error );
  input [31:0] address_bus;
  input [31:0] data_bus;
  input [15:0] dependency_remove;
  output [31:0] read_data_buff;
  output [15:0] instruction_out;
  output [3:0] out_reg;
  input clk, n_rst, read_instruction, valid_data, read_data_enable,
         instruction_buffer_full;
  output add_instruction, read_error, write_error;
  wire   N13, N14, N15, N16, \count[15][3] , \count[15][2] , \count[15][1] ,
         \count[15][0] , \count[14][3] , \count[14][2] , \count[14][1] ,
         \count[14][0] , \count[13][3] , \count[13][2] , \count[13][1] ,
         \count[13][0] , \count[12][3] , \count[12][2] , \count[12][1] ,
         \count[12][0] , \count[11][3] , \count[11][2] , \count[11][1] ,
         \count[11][0] , \count[10][3] , \count[10][2] , \count[10][1] ,
         \count[10][0] , \count[9][3] , \count[9][2] , \count[9][1] ,
         \count[9][0] , \count[8][3] , \count[8][2] , \count[8][1] ,
         \count[8][0] , \count[7][3] , \count[7][2] , \count[7][1] ,
         \count[7][0] , \count[6][3] , \count[6][2] , \count[6][1] ,
         \count[6][0] , \count[5][3] , \count[5][2] , \count[5][1] ,
         \count[5][0] , \count[4][3] , \count[4][2] , \count[4][1] ,
         \count[4][0] , \count[3][3] , \count[3][2] , \count[3][1] ,
         \count[3][0] , \count[2][3] , \count[2][2] , \count[2][1] ,
         \count[2][0] , \count[1][3] , \count[1][2] , \count[1][1] ,
         \count[1][0] , \count[0][3] , \count[0][2] , \count[0][1] ,
         \count[0][0] , fifo_full, prev_fifo, N38, N39, N40, N41, N42, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100;
  wire   [15:0] cnt_up;
  assign out_reg[0] = N13;
  assign N13 = address_bus[0];
  assign out_reg[1] = N14;
  assign N14 = address_bus[1];
  assign out_reg[2] = N15;
  assign N15 = address_bus[2];
  assign out_reg[3] = N16;
  assign N16 = address_bus[3];
  assign instruction_out[15] = address_bus[31];
  assign instruction_out[14] = address_bus[30];
  assign instruction_out[13] = address_bus[29];
  assign instruction_out[12] = address_bus[28];
  assign instruction_out[11] = address_bus[27];
  assign instruction_out[10] = address_bus[26];
  assign instruction_out[9] = address_bus[25];
  assign instruction_out[8] = address_bus[24];
  assign instruction_out[7] = address_bus[23];
  assign instruction_out[6] = address_bus[22];
  assign instruction_out[5] = address_bus[21];
  assign instruction_out[4] = address_bus[20];
  assign instruction_out[3] = address_bus[19];
  assign instruction_out[2] = address_bus[18];
  assign instruction_out[1] = address_bus[17];
  assign instruction_out[0] = address_bus[16];
  assign read_error = N42;

  DFFSR prev_fifo_reg ( .D(fifo_full), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        prev_fifo) );
  AND2X2 U4 ( .A(valid_data), .B(instruction_out[15]), .Y(n13) );
  AND2X2 U5 ( .A(n100), .B(prev_fifo), .Y(n15) );
  AND2X2 U6 ( .A(instruction_out[9]), .B(n26), .Y(n24) );
  AND2X2 U7 ( .A(prev_fifo), .B(fifo_full), .Y(n30) );
  NOR2X1 U17 ( .A(n11), .B(n12), .Y(write_error) );
  NAND3X1 U18 ( .A(instruction_out[13]), .B(fifo_full), .C(n13), .Y(n12) );
  NAND3X1 U19 ( .A(n14), .B(n95), .C(n15), .Y(n11) );
  NOR2X1 U20 ( .A(read_instruction), .B(instruction_out[14]), .Y(n14) );
  NOR2X1 U21 ( .A(n16), .B(n17), .Y(cnt_up[9]) );
  NOR2X1 U22 ( .A(n16), .B(n18), .Y(cnt_up[8]) );
  NOR2X1 U23 ( .A(n19), .B(n20), .Y(cnt_up[7]) );
  NOR2X1 U24 ( .A(n19), .B(n21), .Y(cnt_up[6]) );
  NOR2X1 U25 ( .A(n20), .B(n22), .Y(cnt_up[5]) );
  NOR2X1 U26 ( .A(n21), .B(n22), .Y(cnt_up[4]) );
  NOR2X1 U27 ( .A(n20), .B(n23), .Y(cnt_up[3]) );
  NOR2X1 U28 ( .A(n21), .B(n23), .Y(cnt_up[2]) );
  NOR2X1 U29 ( .A(n16), .B(n20), .Y(cnt_up[1]) );
  NAND2X1 U30 ( .A(instruction_out[8]), .B(n96), .Y(n20) );
  NOR2X1 U31 ( .A(n17), .B(n19), .Y(cnt_up[15]) );
  NOR2X1 U32 ( .A(n18), .B(n19), .Y(cnt_up[14]) );
  NAND2X1 U33 ( .A(instruction_out[10]), .B(n24), .Y(n19) );
  NOR2X1 U34 ( .A(n17), .B(n22), .Y(cnt_up[13]) );
  NOR2X1 U35 ( .A(n18), .B(n22), .Y(cnt_up[12]) );
  NAND2X1 U36 ( .A(instruction_out[10]), .B(n25), .Y(n22) );
  NOR2X1 U37 ( .A(n17), .B(n23), .Y(cnt_up[11]) );
  NAND2X1 U38 ( .A(instruction_out[8]), .B(instruction_out[11]), .Y(n17) );
  NOR2X1 U39 ( .A(n18), .B(n23), .Y(cnt_up[10]) );
  NAND2X1 U40 ( .A(n24), .B(n97), .Y(n23) );
  NAND2X1 U41 ( .A(instruction_out[11]), .B(n98), .Y(n18) );
  NOR2X1 U42 ( .A(n16), .B(n21), .Y(cnt_up[0]) );
  NAND2X1 U43 ( .A(n96), .B(n98), .Y(n21) );
  NAND2X1 U44 ( .A(n25), .B(n97), .Y(n16) );
  NOR2X1 U45 ( .A(n92), .B(instruction_out[9]), .Y(n25) );
  NOR2X1 U46 ( .A(n27), .B(n28), .Y(n26) );
  XOR2X1 U47 ( .A(instruction_out[15]), .B(n29), .Y(n27) );
  NOR2X1 U48 ( .A(instruction_out[13]), .B(instruction_out[14]), .Y(n29) );
  AOI21X1 U49 ( .A(n30), .B(n93), .C(n28), .Y(add_instruction) );
  NAND3X1 U50 ( .A(n32), .B(instruction_out[15]), .C(n33), .Y(n31) );
  NOR2X1 U51 ( .A(n94), .B(n28), .Y(n33) );
  NAND3X1 U52 ( .A(n100), .B(n99), .C(valid_data), .Y(n28) );
  NOR2X1 U53 ( .A(instruction_out[14]), .B(instruction_out[12]), .Y(n32) );
  AOI21X1 U54 ( .A(n34), .B(n35), .C(n99), .Y(N42) );
  NOR2X1 U55 ( .A(N41), .B(N40), .Y(n35) );
  NOR2X1 U56 ( .A(N39), .B(N38), .Y(n34) );
  upDownCounter_15 \genblk1[0].IX  ( .clk(clk), .n_rst(n_rst), .up(cnt_up[0]), 
        .down(dependency_remove[0]), .count_out({\count[0][3] , \count[0][2] , 
        \count[0][1] , \count[0][0] }) );
  upDownCounter_14 \genblk1[1].IX  ( .clk(clk), .n_rst(n_rst), .up(cnt_up[1]), 
        .down(dependency_remove[1]), .count_out({\count[1][3] , \count[1][2] , 
        \count[1][1] , \count[1][0] }) );
  upDownCounter_13 \genblk1[2].IX  ( .clk(clk), .n_rst(n_rst), .up(cnt_up[2]), 
        .down(dependency_remove[2]), .count_out({\count[2][3] , \count[2][2] , 
        \count[2][1] , \count[2][0] }) );
  upDownCounter_12 \genblk1[3].IX  ( .clk(clk), .n_rst(n_rst), .up(cnt_up[3]), 
        .down(dependency_remove[3]), .count_out({\count[3][3] , \count[3][2] , 
        \count[3][1] , \count[3][0] }) );
  upDownCounter_11 \genblk1[4].IX  ( .clk(clk), .n_rst(n_rst), .up(cnt_up[4]), 
        .down(dependency_remove[4]), .count_out({\count[4][3] , \count[4][2] , 
        \count[4][1] , \count[4][0] }) );
  upDownCounter_10 \genblk1[5].IX  ( .clk(clk), .n_rst(n_rst), .up(cnt_up[5]), 
        .down(dependency_remove[5]), .count_out({\count[5][3] , \count[5][2] , 
        \count[5][1] , \count[5][0] }) );
  upDownCounter_9 \genblk1[6].IX  ( .clk(clk), .n_rst(n_rst), .up(cnt_up[6]), 
        .down(dependency_remove[6]), .count_out({\count[6][3] , \count[6][2] , 
        \count[6][1] , \count[6][0] }) );
  upDownCounter_8 \genblk1[7].IX  ( .clk(clk), .n_rst(n_rst), .up(cnt_up[7]), 
        .down(dependency_remove[7]), .count_out({\count[7][3] , \count[7][2] , 
        \count[7][1] , \count[7][0] }) );
  upDownCounter_7 \genblk1[8].IX  ( .clk(clk), .n_rst(n_rst), .up(cnt_up[8]), 
        .down(dependency_remove[8]), .count_out({\count[8][3] , \count[8][2] , 
        \count[8][1] , \count[8][0] }) );
  upDownCounter_6 \genblk1[9].IX  ( .clk(clk), .n_rst(n_rst), .up(cnt_up[9]), 
        .down(dependency_remove[9]), .count_out({\count[9][3] , \count[9][2] , 
        \count[9][1] , \count[9][0] }) );
  upDownCounter_5 \genblk1[10].IX  ( .clk(clk), .n_rst(n_rst), .up(cnt_up[10]), 
        .down(dependency_remove[10]), .count_out({\count[10][3] , 
        \count[10][2] , \count[10][1] , \count[10][0] }) );
  upDownCounter_4 \genblk1[11].IX  ( .clk(clk), .n_rst(n_rst), .up(cnt_up[11]), 
        .down(dependency_remove[11]), .count_out({\count[11][3] , 
        \count[11][2] , \count[11][1] , \count[11][0] }) );
  upDownCounter_3 \genblk1[12].IX  ( .clk(clk), .n_rst(n_rst), .up(cnt_up[12]), 
        .down(dependency_remove[12]), .count_out({\count[12][3] , 
        \count[12][2] , \count[12][1] , \count[12][0] }) );
  upDownCounter_2 \genblk1[13].IX  ( .clk(clk), .n_rst(n_rst), .up(cnt_up[13]), 
        .down(dependency_remove[13]), .count_out({\count[13][3] , 
        \count[13][2] , \count[13][1] , \count[13][0] }) );
  upDownCounter_1 \genblk1[14].IX  ( .clk(clk), .n_rst(n_rst), .up(cnt_up[14]), 
        .down(dependency_remove[14]), .count_out({\count[14][3] , 
        \count[14][2] , \count[14][1] , \count[14][0] }) );
  upDownCounter_0 \genblk1[15].IX  ( .clk(clk), .n_rst(n_rst), .up(cnt_up[15]), 
        .down(dependency_remove[15]), .count_out({\count[15][3] , 
        \count[15][2] , \count[15][1] , \count[15][0] }) );
  flex_fifo_WIDTH32_DEPTH4_BITS_WIDTH5_BITS_DEPTH2 Data_buffer ( .clk(clk), 
        .n_rst(n_rst), .r_enable(read_data_enable), .w_enable(n93), .w_data(
        data_bus), .r_data(read_data_buff), .full(fifo_full) );
  MUX2X1 U57 ( .B(n37), .A(n38), .S(N14), .Y(n36) );
  MUX2X1 U58 ( .B(n40), .A(n41), .S(N14), .Y(n39) );
  MUX2X1 U59 ( .B(n43), .A(n44), .S(N14), .Y(n42) );
  MUX2X1 U60 ( .B(n46), .A(n47), .S(N14), .Y(n45) );
  MUX2X1 U61 ( .B(n48), .A(n49), .S(N16), .Y(N41) );
  MUX2X1 U62 ( .B(n51), .A(n52), .S(N14), .Y(n50) );
  MUX2X1 U63 ( .B(n54), .A(n55), .S(N14), .Y(n53) );
  MUX2X1 U64 ( .B(n57), .A(n58), .S(N14), .Y(n56) );
  MUX2X1 U65 ( .B(n60), .A(n61), .S(N14), .Y(n59) );
  MUX2X1 U66 ( .B(n62), .A(n63), .S(N16), .Y(N40) );
  MUX2X1 U67 ( .B(n65), .A(n66), .S(N14), .Y(n64) );
  MUX2X1 U68 ( .B(n68), .A(n69), .S(N14), .Y(n67) );
  MUX2X1 U69 ( .B(n71), .A(n72), .S(N14), .Y(n70) );
  MUX2X1 U70 ( .B(n74), .A(n75), .S(N14), .Y(n73) );
  MUX2X1 U71 ( .B(n76), .A(n77), .S(N16), .Y(N39) );
  MUX2X1 U72 ( .B(n79), .A(n80), .S(N14), .Y(n78) );
  MUX2X1 U73 ( .B(n82), .A(n83), .S(N14), .Y(n81) );
  MUX2X1 U74 ( .B(n85), .A(n86), .S(N14), .Y(n84) );
  MUX2X1 U75 ( .B(n88), .A(n89), .S(N14), .Y(n87) );
  MUX2X1 U76 ( .B(n90), .A(n91), .S(N16), .Y(N38) );
  MUX2X1 U77 ( .B(\count[14][0] ), .A(\count[15][0] ), .S(N13), .Y(n38) );
  MUX2X1 U78 ( .B(\count[12][0] ), .A(\count[13][0] ), .S(N13), .Y(n37) );
  MUX2X1 U79 ( .B(\count[10][0] ), .A(\count[11][0] ), .S(N13), .Y(n41) );
  MUX2X1 U80 ( .B(\count[8][0] ), .A(\count[9][0] ), .S(N13), .Y(n40) );
  MUX2X1 U81 ( .B(n39), .A(n36), .S(N15), .Y(n49) );
  MUX2X1 U82 ( .B(\count[6][0] ), .A(\count[7][0] ), .S(N13), .Y(n44) );
  MUX2X1 U83 ( .B(\count[4][0] ), .A(\count[5][0] ), .S(N13), .Y(n43) );
  MUX2X1 U84 ( .B(\count[2][0] ), .A(\count[3][0] ), .S(N13), .Y(n47) );
  MUX2X1 U85 ( .B(\count[0][0] ), .A(\count[1][0] ), .S(N13), .Y(n46) );
  MUX2X1 U86 ( .B(n45), .A(n42), .S(N15), .Y(n48) );
  MUX2X1 U87 ( .B(\count[14][1] ), .A(\count[15][1] ), .S(N13), .Y(n52) );
  MUX2X1 U88 ( .B(\count[12][1] ), .A(\count[13][1] ), .S(N13), .Y(n51) );
  MUX2X1 U89 ( .B(\count[10][1] ), .A(\count[11][1] ), .S(N13), .Y(n55) );
  MUX2X1 U90 ( .B(\count[8][1] ), .A(\count[9][1] ), .S(N13), .Y(n54) );
  MUX2X1 U91 ( .B(n53), .A(n50), .S(N15), .Y(n63) );
  MUX2X1 U92 ( .B(\count[6][1] ), .A(\count[7][1] ), .S(N13), .Y(n58) );
  MUX2X1 U93 ( .B(\count[4][1] ), .A(\count[5][1] ), .S(N13), .Y(n57) );
  MUX2X1 U94 ( .B(\count[2][1] ), .A(\count[3][1] ), .S(N13), .Y(n61) );
  MUX2X1 U95 ( .B(\count[0][1] ), .A(\count[1][1] ), .S(N13), .Y(n60) );
  MUX2X1 U96 ( .B(n59), .A(n56), .S(N15), .Y(n62) );
  MUX2X1 U97 ( .B(\count[14][2] ), .A(\count[15][2] ), .S(N13), .Y(n66) );
  MUX2X1 U98 ( .B(\count[12][2] ), .A(\count[13][2] ), .S(N13), .Y(n65) );
  MUX2X1 U99 ( .B(\count[10][2] ), .A(\count[11][2] ), .S(N13), .Y(n69) );
  MUX2X1 U100 ( .B(\count[8][2] ), .A(\count[9][2] ), .S(N13), .Y(n68) );
  MUX2X1 U101 ( .B(n67), .A(n64), .S(N15), .Y(n77) );
  MUX2X1 U102 ( .B(\count[6][2] ), .A(\count[7][2] ), .S(N13), .Y(n72) );
  MUX2X1 U103 ( .B(\count[4][2] ), .A(\count[5][2] ), .S(N13), .Y(n71) );
  MUX2X1 U104 ( .B(\count[2][2] ), .A(\count[3][2] ), .S(N13), .Y(n75) );
  MUX2X1 U105 ( .B(\count[0][2] ), .A(\count[1][2] ), .S(N13), .Y(n74) );
  MUX2X1 U106 ( .B(n73), .A(n70), .S(N15), .Y(n76) );
  MUX2X1 U107 ( .B(\count[14][3] ), .A(\count[15][3] ), .S(N13), .Y(n80) );
  MUX2X1 U108 ( .B(\count[12][3] ), .A(\count[13][3] ), .S(N13), .Y(n79) );
  MUX2X1 U109 ( .B(\count[10][3] ), .A(\count[11][3] ), .S(N13), .Y(n83) );
  MUX2X1 U110 ( .B(\count[8][3] ), .A(\count[9][3] ), .S(N13), .Y(n82) );
  MUX2X1 U111 ( .B(n81), .A(n78), .S(N15), .Y(n91) );
  MUX2X1 U112 ( .B(\count[6][3] ), .A(\count[7][3] ), .S(N13), .Y(n86) );
  MUX2X1 U113 ( .B(\count[4][3] ), .A(\count[5][3] ), .S(N13), .Y(n85) );
  MUX2X1 U114 ( .B(\count[2][3] ), .A(\count[3][3] ), .S(N13), .Y(n89) );
  MUX2X1 U115 ( .B(\count[0][3] ), .A(\count[1][3] ), .S(N13), .Y(n88) );
  MUX2X1 U116 ( .B(n87), .A(n84), .S(N15), .Y(n90) );
  INVX2 U117 ( .A(n26), .Y(n92) );
  INVX2 U118 ( .A(n31), .Y(n93) );
  INVX2 U119 ( .A(instruction_out[13]), .Y(n94) );
  INVX2 U120 ( .A(instruction_out[12]), .Y(n95) );
  INVX2 U121 ( .A(instruction_out[11]), .Y(n96) );
  INVX2 U122 ( .A(instruction_out[10]), .Y(n97) );
  INVX2 U123 ( .A(instruction_out[8]), .Y(n98) );
  INVX2 U124 ( .A(read_instruction), .Y(n99) );
  INVX2 U125 ( .A(instruction_buffer_full), .Y(n100) );
endmodule

