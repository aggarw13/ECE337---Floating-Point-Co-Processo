
module flex_indexer_NUM_CNT_BITS3_1 ( clk, n_rst, clear, count_enable, 
        rollover_val, count_out, rollover_flag );
  input [2:0] rollover_val;
  output [2:0] count_out;
  input clk, n_rst, clear, count_enable;
  output rollover_flag;
  wire   n27, n28, n2, n3, n4, n8, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26;
  wire   [2:0] nxt_count;
  assign rollover_flag = 1'b0;

  DFFSR \count_out_reg[0]  ( .D(nxt_count[0]), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(n28) );
  DFFSR \count_out_reg[2]  ( .D(nxt_count[2]), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(n27) );
  DFFSR \count_out_reg[1]  ( .D(nxt_count[1]), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(count_out[1]) );
  INVX2 U7 ( .A(n2), .Y(n3) );
  BUFX4 U8 ( .A(n28), .Y(count_out[0]) );
  INVX1 U9 ( .A(count_out[1]), .Y(n2) );
  INVX1 U10 ( .A(n20), .Y(n4) );
  INVX1 U11 ( .A(count_out[0]), .Y(n20) );
  INVX2 U12 ( .A(n27), .Y(n8) );
  INVX4 U13 ( .A(n8), .Y(count_out[2]) );
  BUFX2 U14 ( .A(n3), .Y(n10) );
  INVX2 U15 ( .A(clear), .Y(n17) );
  INVX2 U16 ( .A(count_out[2]), .Y(n22) );
  XOR2X1 U17 ( .A(n22), .B(rollover_val[2]), .Y(n13) );
  XOR2X1 U18 ( .A(n20), .B(rollover_val[0]), .Y(n12) );
  XNOR2X1 U19 ( .A(n3), .B(rollover_val[1]), .Y(n11) );
  NAND3X1 U20 ( .A(n13), .B(n12), .C(n11), .Y(n14) );
  NAND3X1 U21 ( .A(n17), .B(n14), .C(count_enable), .Y(n26) );
  INVX2 U22 ( .A(n26), .Y(n15) );
  NAND2X1 U23 ( .A(n15), .B(n4), .Y(n19) );
  INVX2 U24 ( .A(count_enable), .Y(n16) );
  NAND2X1 U25 ( .A(n17), .B(n16), .Y(n25) );
  OAI21X1 U26 ( .A(n4), .B(n26), .C(n25), .Y(n18) );
  INVX2 U27 ( .A(n18), .Y(n23) );
  MUX2X1 U28 ( .B(n19), .A(n23), .S(n10), .Y(nxt_count[1]) );
  NOR2X1 U29 ( .A(count_out[2]), .B(n20), .Y(n21) );
  MUX2X1 U30 ( .B(count_out[2]), .A(n21), .S(n10), .Y(n24) );
  OAI22X1 U31 ( .A(n24), .B(n26), .C(n23), .D(n22), .Y(nxt_count[2]) );
  MUX2X1 U32 ( .B(n26), .A(n25), .S(n4), .Y(nxt_count[0]) );
endmodule


module flex_indexer_NUM_CNT_BITS3_0 ( clk, n_rst, clear, count_enable, 
        rollover_val, count_out, rollover_flag );
  input [2:0] rollover_val;
  output [2:0] count_out;
  input clk, n_rst, clear, count_enable;
  output rollover_flag;
  wire   n29, n30, n31, n1, n2, n4, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25;
  wire   [2:0] nxt_count;
  assign rollover_flag = 1'b0;

  DFFSR \count_out_reg[0]  ( .D(nxt_count[0]), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(n31) );
  DFFSR \count_out_reg[2]  ( .D(nxt_count[2]), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(n29) );
  DFFSR \count_out_reg[1]  ( .D(nxt_count[1]), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(n30) );
  BUFX2 U7 ( .A(count_out[1]), .Y(n1) );
  INVX4 U8 ( .A(n31), .Y(n10) );
  BUFX2 U9 ( .A(n1), .Y(n2) );
  BUFX4 U10 ( .A(n30), .Y(count_out[1]) );
  INVX2 U11 ( .A(n29), .Y(n4) );
  INVX8 U12 ( .A(n4), .Y(count_out[2]) );
  INVX8 U13 ( .A(n10), .Y(count_out[0]) );
  INVX2 U14 ( .A(count_out[2]), .Y(n21) );
  XOR2X1 U15 ( .A(n21), .B(rollover_val[2]), .Y(n13) );
  XOR2X1 U16 ( .A(n10), .B(rollover_val[0]), .Y(n12) );
  XNOR2X1 U17 ( .A(n1), .B(rollover_val[1]), .Y(n11) );
  NAND3X1 U18 ( .A(n13), .B(n12), .C(n11), .Y(n16) );
  INVX2 U19 ( .A(clear), .Y(n17) );
  NAND3X1 U20 ( .A(n16), .B(n17), .C(count_enable), .Y(n25) );
  INVX2 U21 ( .A(n25), .Y(n14) );
  NAND2X1 U22 ( .A(n14), .B(count_out[0]), .Y(n19) );
  INVX2 U23 ( .A(count_enable), .Y(n15) );
  NAND2X1 U24 ( .A(n17), .B(n15), .Y(n24) );
  NAND3X1 U25 ( .A(n17), .B(n10), .C(n16), .Y(n18) );
  AND2X2 U26 ( .A(n24), .B(n18), .Y(n22) );
  MUX2X1 U27 ( .B(n19), .A(n22), .S(n2), .Y(nxt_count[1]) );
  NOR2X1 U28 ( .A(count_out[2]), .B(n10), .Y(n20) );
  MUX2X1 U29 ( .B(count_out[2]), .A(n20), .S(n2), .Y(n23) );
  OAI22X1 U30 ( .A(n23), .B(n25), .C(n22), .D(n21), .Y(nxt_count[2]) );
  MUX2X1 U31 ( .B(n25), .A(n24), .S(count_out[0]), .Y(nxt_count[0]) );
endmodule


module flex_fifo ( clk, n_rst, r_enable, w_enable, w_data, r_data, full, empty
 );
  input [7:0] w_data;
  output [7:0] r_data;
  input clk, n_rst, r_enable, w_enable;
  output full, empty;
  wire   N8, N9, N10, _1_net_, \data[7][7] , \data[7][6] , \data[7][5] ,
         \data[7][4] , \data[7][3] , \data[7][2] , \data[7][1] , \data[7][0] ,
         \data[6][7] , \data[6][6] , \data[6][5] , \data[6][4] , \data[6][3] ,
         \data[6][2] , \data[6][1] , \data[6][0] , \data[5][7] , \data[5][6] ,
         \data[5][5] , \data[5][4] , \data[5][3] , \data[5][2] , \data[5][1] ,
         \data[5][0] , \data[4][7] , \data[4][6] , \data[4][5] , \data[4][4] ,
         \data[4][3] , \data[4][2] , \data[4][1] , \data[4][0] , \data[3][7] ,
         \data[3][6] , \data[3][5] , \data[3][4] , \data[3][3] , \data[3][2] ,
         \data[3][1] , \data[3][0] , \data[2][7] , \data[2][6] , \data[2][5] ,
         \data[2][4] , \data[2][3] , \data[2][2] , \data[2][1] , \data[2][0] ,
         \data[1][7] , \data[1][6] , \data[1][5] , \data[1][4] , \data[1][3] ,
         \data[1][2] , \data[1][1] , \data[1][0] , \data[0][7] , \data[0][6] ,
         \data[0][5] , \data[0][4] , \data[0][3] , \data[0][2] , \data[0][1] ,
         \data[0][0] , \nxt_data[7][7] , \nxt_data[7][6] , \nxt_data[7][5] ,
         \nxt_data[7][4] , \nxt_data[7][3] , \nxt_data[7][2] ,
         \nxt_data[7][1] , \nxt_data[7][0] , \nxt_data[6][7] ,
         \nxt_data[6][6] , \nxt_data[6][5] , \nxt_data[6][4] ,
         \nxt_data[6][3] , \nxt_data[6][2] , \nxt_data[6][1] ,
         \nxt_data[6][0] , \nxt_data[5][7] , \nxt_data[5][6] ,
         \nxt_data[5][5] , \nxt_data[5][4] , \nxt_data[5][3] ,
         \nxt_data[5][2] , \nxt_data[5][1] , \nxt_data[5][0] ,
         \nxt_data[4][7] , \nxt_data[4][6] , \nxt_data[4][5] ,
         \nxt_data[4][4] , \nxt_data[4][3] , \nxt_data[4][2] ,
         \nxt_data[4][1] , \nxt_data[4][0] , \nxt_data[3][7] ,
         \nxt_data[3][6] , \nxt_data[3][5] , \nxt_data[3][4] ,
         \nxt_data[3][3] , \nxt_data[3][2] , \nxt_data[3][1] ,
         \nxt_data[3][0] , \nxt_data[2][7] , \nxt_data[2][6] ,
         \nxt_data[2][5] , \nxt_data[2][4] , \nxt_data[2][3] ,
         \nxt_data[2][2] , \nxt_data[2][1] , \nxt_data[2][0] ,
         \nxt_data[1][7] , \nxt_data[1][6] , \nxt_data[1][5] ,
         \nxt_data[1][4] , \nxt_data[1][3] , \nxt_data[1][2] ,
         \nxt_data[1][1] , \nxt_data[1][0] , \nxt_data[0][7] ,
         \nxt_data[0][6] , \nxt_data[0][5] , \nxt_data[0][4] ,
         \nxt_data[0][3] , \nxt_data[0][2] , \nxt_data[0][1] ,
         \nxt_data[0][0] , n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385;
  wire   [2:0] w_pointer;

  DFFSR \data_reg[7][7]  ( .D(\nxt_data[7][7] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[7][7] ) );
  DFFSR \data_reg[7][6]  ( .D(\nxt_data[7][6] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[7][6] ) );
  DFFSR \data_reg[7][5]  ( .D(\nxt_data[7][5] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[7][5] ) );
  DFFSR \data_reg[7][4]  ( .D(\nxt_data[7][4] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[7][4] ) );
  DFFSR \data_reg[7][3]  ( .D(\nxt_data[7][3] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[7][3] ) );
  DFFSR \data_reg[7][2]  ( .D(\nxt_data[7][2] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[7][2] ) );
  DFFSR \data_reg[7][1]  ( .D(\nxt_data[7][1] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[7][1] ) );
  DFFSR \data_reg[7][0]  ( .D(\nxt_data[7][0] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[7][0] ) );
  DFFSR \data_reg[6][7]  ( .D(\nxt_data[6][7] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[6][7] ) );
  DFFSR \data_reg[6][6]  ( .D(\nxt_data[6][6] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[6][6] ) );
  DFFSR \data_reg[6][5]  ( .D(\nxt_data[6][5] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[6][5] ) );
  DFFSR \data_reg[6][4]  ( .D(\nxt_data[6][4] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[6][4] ) );
  DFFSR \data_reg[6][3]  ( .D(\nxt_data[6][3] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[6][3] ) );
  DFFSR \data_reg[6][2]  ( .D(\nxt_data[6][2] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[6][2] ) );
  DFFSR \data_reg[6][1]  ( .D(\nxt_data[6][1] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[6][1] ) );
  DFFSR \data_reg[6][0]  ( .D(\nxt_data[6][0] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[6][0] ) );
  DFFSR \data_reg[5][7]  ( .D(\nxt_data[5][7] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[5][7] ) );
  DFFSR \data_reg[5][6]  ( .D(\nxt_data[5][6] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[5][6] ) );
  DFFSR \data_reg[5][5]  ( .D(\nxt_data[5][5] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[5][5] ) );
  DFFSR \data_reg[5][4]  ( .D(\nxt_data[5][4] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[5][4] ) );
  DFFSR \data_reg[5][3]  ( .D(\nxt_data[5][3] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[5][3] ) );
  DFFSR \data_reg[5][2]  ( .D(\nxt_data[5][2] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[5][2] ) );
  DFFSR \data_reg[5][1]  ( .D(\nxt_data[5][1] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[5][1] ) );
  DFFSR \data_reg[5][0]  ( .D(\nxt_data[5][0] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[5][0] ) );
  DFFSR \data_reg[4][7]  ( .D(\nxt_data[4][7] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[4][7] ) );
  DFFSR \data_reg[4][6]  ( .D(\nxt_data[4][6] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[4][6] ) );
  DFFSR \data_reg[4][5]  ( .D(\nxt_data[4][5] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[4][5] ) );
  DFFSR \data_reg[4][4]  ( .D(\nxt_data[4][4] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[4][4] ) );
  DFFSR \data_reg[4][3]  ( .D(\nxt_data[4][3] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[4][3] ) );
  DFFSR \data_reg[4][2]  ( .D(\nxt_data[4][2] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[4][2] ) );
  DFFSR \data_reg[4][1]  ( .D(\nxt_data[4][1] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[4][1] ) );
  DFFSR \data_reg[4][0]  ( .D(\nxt_data[4][0] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[4][0] ) );
  DFFSR \data_reg[3][7]  ( .D(\nxt_data[3][7] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[3][7] ) );
  DFFSR \data_reg[3][6]  ( .D(\nxt_data[3][6] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[3][6] ) );
  DFFSR \data_reg[3][5]  ( .D(\nxt_data[3][5] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[3][5] ) );
  DFFSR \data_reg[3][4]  ( .D(\nxt_data[3][4] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[3][4] ) );
  DFFSR \data_reg[3][3]  ( .D(\nxt_data[3][3] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[3][3] ) );
  DFFSR \data_reg[3][2]  ( .D(\nxt_data[3][2] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[3][2] ) );
  DFFSR \data_reg[3][1]  ( .D(\nxt_data[3][1] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[3][1] ) );
  DFFSR \data_reg[3][0]  ( .D(\nxt_data[3][0] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[3][0] ) );
  DFFSR \data_reg[2][7]  ( .D(\nxt_data[2][7] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[2][7] ) );
  DFFSR \data_reg[2][6]  ( .D(\nxt_data[2][6] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[2][6] ) );
  DFFSR \data_reg[2][5]  ( .D(\nxt_data[2][5] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[2][5] ) );
  DFFSR \data_reg[2][4]  ( .D(\nxt_data[2][4] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[2][4] ) );
  DFFSR \data_reg[2][3]  ( .D(\nxt_data[2][3] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[2][3] ) );
  DFFSR \data_reg[2][2]  ( .D(\nxt_data[2][2] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[2][2] ) );
  DFFSR \data_reg[2][1]  ( .D(\nxt_data[2][1] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[2][1] ) );
  DFFSR \data_reg[2][0]  ( .D(\nxt_data[2][0] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[2][0] ) );
  DFFSR \data_reg[1][7]  ( .D(\nxt_data[1][7] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[1][7] ) );
  DFFSR \data_reg[1][6]  ( .D(\nxt_data[1][6] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[1][6] ) );
  DFFSR \data_reg[1][5]  ( .D(\nxt_data[1][5] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[1][5] ) );
  DFFSR \data_reg[1][4]  ( .D(\nxt_data[1][4] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[1][4] ) );
  DFFSR \data_reg[1][3]  ( .D(\nxt_data[1][3] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[1][3] ) );
  DFFSR \data_reg[1][2]  ( .D(\nxt_data[1][2] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[1][2] ) );
  DFFSR \data_reg[1][1]  ( .D(\nxt_data[1][1] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[1][1] ) );
  DFFSR \data_reg[1][0]  ( .D(\nxt_data[1][0] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[1][0] ) );
  DFFSR \data_reg[0][7]  ( .D(\nxt_data[0][7] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[0][7] ) );
  DFFSR \data_reg[0][6]  ( .D(\nxt_data[0][6] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[0][6] ) );
  DFFSR \data_reg[0][5]  ( .D(\nxt_data[0][5] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[0][5] ) );
  DFFSR \data_reg[0][4]  ( .D(\nxt_data[0][4] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[0][4] ) );
  DFFSR \data_reg[0][3]  ( .D(\nxt_data[0][3] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[0][3] ) );
  DFFSR \data_reg[0][2]  ( .D(\nxt_data[0][2] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[0][2] ) );
  DFFSR \data_reg[0][1]  ( .D(\nxt_data[0][1] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[0][1] ) );
  DFFSR \data_reg[0][0]  ( .D(\nxt_data[0][0] ), .CLK(clk), .R(n_rst), .S(1'b1), .Q(\data[0][0] ) );
  flex_indexer_NUM_CNT_BITS3_1 Write_pointer ( .clk(clk), .n_rst(n_rst), 
        .clear(1'b0), .count_enable(w_enable), .rollover_val({1'b1, 1'b1, 1'b1}), .count_out(w_pointer) );
  flex_indexer_NUM_CNT_BITS3_0 Read_pointer ( .clk(clk), .n_rst(n_rst), 
        .clear(1'b0), .count_enable(_1_net_), .rollover_val({1'b1, 1'b1, 1'b1}), .count_out({N10, N9, N8}) );
  INVX1 U235 ( .A(n330), .Y(n178) );
  INVX2 U236 ( .A(n330), .Y(n334) );
  AND2X2 U237 ( .A(w_enable), .B(n280), .Y(n179) );
  INVX2 U238 ( .A(w_pointer[2]), .Y(n280) );
  INVX1 U239 ( .A(n273), .Y(empty) );
  INVX1 U240 ( .A(n356), .Y(n180) );
  INVX1 U241 ( .A(n348), .Y(n181) );
  INVX1 U242 ( .A(n348), .Y(n352) );
  INVX1 U243 ( .A(n348), .Y(n182) );
  INVX1 U244 ( .A(n348), .Y(n183) );
  INVX2 U245 ( .A(n186), .Y(n257) );
  INVX2 U246 ( .A(n336), .Y(n186) );
  MUX2X1 U247 ( .B(n342), .A(n372), .S(n184), .Y(\nxt_data[5][1] ) );
  INVX1 U248 ( .A(n340), .Y(n184) );
  BUFX2 U249 ( .A(n363), .Y(n185) );
  BUFX2 U250 ( .A(n363), .Y(n187) );
  MUX2X1 U251 ( .B(n341), .A(n370), .S(n344), .Y(\nxt_data[5][0] ) );
  NAND2X1 U252 ( .A(n286), .B(n329), .Y(n188) );
  INVX2 U253 ( .A(w_pointer[1]), .Y(n336) );
  AND2X2 U254 ( .A(n279), .B(n278), .Y(n189) );
  BUFX4 U255 ( .A(w_pointer[0]), .Y(n254) );
  INVX2 U256 ( .A(n249), .Y(n250) );
  INVX2 U257 ( .A(n249), .Y(n251) );
  INVX2 U258 ( .A(n253), .Y(n252) );
  INVX1 U259 ( .A(N8), .Y(n249) );
  AND2X2 U260 ( .A(n258), .B(n192), .Y(n190) );
  AND2X2 U261 ( .A(n179), .B(n369), .Y(n191) );
  MUX2X1 U262 ( .B(n370), .A(n357), .S(n185), .Y(\nxt_data[6][0] ) );
  MUX2X1 U263 ( .B(n372), .A(n358), .S(n187), .Y(\nxt_data[6][1] ) );
  MUX2X1 U264 ( .B(n382), .A(n366), .S(n185), .Y(\nxt_data[6][6] ) );
  MUX2X1 U265 ( .B(n384), .A(n368), .S(n187), .Y(\nxt_data[6][7] ) );
  MUX2X1 U266 ( .B(n374), .A(n326), .S(n188), .Y(\nxt_data[4][2] ) );
  MUX2X1 U267 ( .B(n376), .A(n328), .S(n188), .Y(\nxt_data[4][3] ) );
  AND2X2 U268 ( .A(w_enable), .B(w_pointer[2]), .Y(n192) );
  MUX2X1 U269 ( .B(n194), .A(n195), .S(n252), .Y(n193) );
  MUX2X1 U270 ( .B(n197), .A(n198), .S(n252), .Y(n196) );
  MUX2X1 U271 ( .B(n200), .A(n201), .S(n252), .Y(n199) );
  MUX2X1 U272 ( .B(n203), .A(n204), .S(n252), .Y(n202) );
  MUX2X1 U273 ( .B(n206), .A(n207), .S(n252), .Y(n205) );
  MUX2X1 U274 ( .B(n209), .A(n210), .S(n252), .Y(n208) );
  MUX2X1 U275 ( .B(n212), .A(n213), .S(n252), .Y(n211) );
  MUX2X1 U276 ( .B(n215), .A(n216), .S(n252), .Y(n214) );
  MUX2X1 U277 ( .B(n218), .A(n219), .S(n252), .Y(n217) );
  MUX2X1 U278 ( .B(n221), .A(n222), .S(n252), .Y(n220) );
  MUX2X1 U279 ( .B(n224), .A(n225), .S(n252), .Y(n223) );
  MUX2X1 U280 ( .B(n227), .A(n228), .S(n252), .Y(n226) );
  MUX2X1 U281 ( .B(n230), .A(n231), .S(n252), .Y(n229) );
  MUX2X1 U282 ( .B(n233), .A(n234), .S(n252), .Y(n232) );
  MUX2X1 U283 ( .B(n236), .A(n237), .S(n252), .Y(n235) );
  MUX2X1 U284 ( .B(n239), .A(n240), .S(n252), .Y(n238) );
  MUX2X1 U285 ( .B(\data[6][0] ), .A(\data[7][0] ), .S(n250), .Y(n195) );
  MUX2X1 U286 ( .B(\data[4][0] ), .A(\data[5][0] ), .S(n251), .Y(n194) );
  MUX2X1 U287 ( .B(\data[2][0] ), .A(\data[3][0] ), .S(n250), .Y(n198) );
  MUX2X1 U288 ( .B(\data[0][0] ), .A(\data[1][0] ), .S(n251), .Y(n197) );
  MUX2X1 U289 ( .B(n196), .A(n193), .S(N10), .Y(n241) );
  MUX2X1 U290 ( .B(\data[6][1] ), .A(\data[7][1] ), .S(n250), .Y(n201) );
  MUX2X1 U291 ( .B(\data[4][1] ), .A(\data[5][1] ), .S(n251), .Y(n200) );
  MUX2X1 U292 ( .B(\data[2][1] ), .A(\data[3][1] ), .S(n250), .Y(n204) );
  MUX2X1 U293 ( .B(\data[0][1] ), .A(\data[1][1] ), .S(n250), .Y(n203) );
  MUX2X1 U294 ( .B(n202), .A(n199), .S(N10), .Y(n242) );
  MUX2X1 U295 ( .B(\data[6][2] ), .A(\data[7][2] ), .S(n250), .Y(n207) );
  MUX2X1 U296 ( .B(\data[4][2] ), .A(\data[5][2] ), .S(n250), .Y(n206) );
  MUX2X1 U297 ( .B(\data[2][2] ), .A(\data[3][2] ), .S(n250), .Y(n210) );
  MUX2X1 U298 ( .B(\data[0][2] ), .A(\data[1][2] ), .S(n250), .Y(n209) );
  MUX2X1 U299 ( .B(n208), .A(n205), .S(N10), .Y(n243) );
  MUX2X1 U300 ( .B(\data[6][3] ), .A(\data[7][3] ), .S(n250), .Y(n213) );
  MUX2X1 U301 ( .B(\data[4][3] ), .A(\data[5][3] ), .S(n250), .Y(n212) );
  MUX2X1 U302 ( .B(\data[2][3] ), .A(\data[3][3] ), .S(n250), .Y(n216) );
  MUX2X1 U303 ( .B(\data[0][3] ), .A(\data[1][3] ), .S(n250), .Y(n215) );
  MUX2X1 U304 ( .B(n214), .A(n211), .S(N10), .Y(n244) );
  MUX2X1 U305 ( .B(\data[6][4] ), .A(\data[7][4] ), .S(n250), .Y(n219) );
  MUX2X1 U306 ( .B(\data[4][4] ), .A(\data[5][4] ), .S(n250), .Y(n218) );
  MUX2X1 U307 ( .B(\data[2][4] ), .A(\data[3][4] ), .S(n250), .Y(n222) );
  MUX2X1 U308 ( .B(\data[0][4] ), .A(\data[1][4] ), .S(n251), .Y(n221) );
  MUX2X1 U309 ( .B(n220), .A(n217), .S(N10), .Y(n245) );
  MUX2X1 U310 ( .B(\data[6][5] ), .A(\data[7][5] ), .S(n251), .Y(n225) );
  MUX2X1 U311 ( .B(\data[4][5] ), .A(\data[5][5] ), .S(n251), .Y(n224) );
  MUX2X1 U312 ( .B(\data[2][5] ), .A(\data[3][5] ), .S(n251), .Y(n228) );
  MUX2X1 U313 ( .B(\data[0][5] ), .A(\data[1][5] ), .S(n251), .Y(n227) );
  MUX2X1 U314 ( .B(n226), .A(n223), .S(N10), .Y(n246) );
  MUX2X1 U315 ( .B(\data[6][6] ), .A(\data[7][6] ), .S(n251), .Y(n231) );
  MUX2X1 U316 ( .B(\data[4][6] ), .A(\data[5][6] ), .S(n251), .Y(n230) );
  MUX2X1 U317 ( .B(\data[2][6] ), .A(\data[3][6] ), .S(n251), .Y(n234) );
  MUX2X1 U318 ( .B(\data[0][6] ), .A(\data[1][6] ), .S(n251), .Y(n233) );
  MUX2X1 U319 ( .B(n232), .A(n229), .S(N10), .Y(n247) );
  MUX2X1 U320 ( .B(\data[6][7] ), .A(\data[7][7] ), .S(n251), .Y(n237) );
  MUX2X1 U321 ( .B(\data[4][7] ), .A(\data[5][7] ), .S(n251), .Y(n236) );
  MUX2X1 U322 ( .B(\data[2][7] ), .A(\data[3][7] ), .S(n251), .Y(n240) );
  MUX2X1 U323 ( .B(\data[0][7] ), .A(\data[1][7] ), .S(n251), .Y(n239) );
  MUX2X1 U324 ( .B(n238), .A(n235), .S(N10), .Y(n248) );
  INVX2 U325 ( .A(n241), .Y(r_data[0]) );
  INVX2 U326 ( .A(n242), .Y(r_data[1]) );
  INVX2 U327 ( .A(n243), .Y(r_data[2]) );
  INVX2 U328 ( .A(n244), .Y(r_data[3]) );
  INVX2 U329 ( .A(n245), .Y(r_data[4]) );
  INVX2 U330 ( .A(n246), .Y(r_data[5]) );
  INVX2 U331 ( .A(n247), .Y(r_data[6]) );
  INVX2 U332 ( .A(n248), .Y(r_data[7]) );
  INVX1 U333 ( .A(N9), .Y(n253) );
  INVX2 U334 ( .A(n257), .Y(n255) );
  BUFX2 U335 ( .A(n254), .Y(n256) );
  INVX1 U336 ( .A(n276), .Y(n258) );
  AOI22X1 U337 ( .A(n276), .B(n277), .C(n369), .D(n275), .Y(n259) );
  INVX1 U338 ( .A(n261), .Y(n260) );
  BUFX2 U339 ( .A(w_pointer[1]), .Y(n261) );
  AND2X2 U340 ( .A(n287), .B(n286), .Y(n262) );
  AND2X2 U341 ( .A(n287), .B(n286), .Y(n263) );
  AND2X2 U342 ( .A(n191), .B(n317), .Y(n264) );
  AND2X2 U343 ( .A(n308), .B(n307), .Y(n265) );
  AND2X2 U344 ( .A(n191), .B(n317), .Y(n266) );
  AND2X2 U345 ( .A(n297), .B(n307), .Y(n267) );
  AND2X2 U346 ( .A(n308), .B(n317), .Y(n268) );
  AND2X2 U347 ( .A(n297), .B(n307), .Y(n269) );
  INVX1 U348 ( .A(n346), .Y(full) );
  XOR2X1 U349 ( .A(n280), .B(N10), .Y(n272) );
  XOR2X1 U350 ( .A(n257), .B(N9), .Y(n271) );
  INVX2 U351 ( .A(w_pointer[0]), .Y(n354) );
  XOR2X1 U352 ( .A(n354), .B(N8), .Y(n270) );
  NAND3X1 U353 ( .A(n272), .B(n271), .C(n270), .Y(n273) );
  AND2X2 U354 ( .A(r_enable), .B(n273), .Y(_1_net_) );
  XOR2X1 U355 ( .A(N10), .B(w_pointer[2]), .Y(n277) );
  NAND2X1 U356 ( .A(w_pointer[0]), .B(n261), .Y(n276) );
  NAND2X1 U357 ( .A(w_pointer[0]), .B(n261), .Y(n274) );
  INVX2 U358 ( .A(n274), .Y(n369) );
  NAND2X1 U359 ( .A(N10), .B(n280), .Y(n275) );
  AOI22X1 U360 ( .A(n277), .B(n276), .C(n369), .D(n275), .Y(n339) );
  FAX1 U361 ( .A(w_pointer[0]), .B(N9), .C(n336), .YS(n279) );
  XOR2X1 U362 ( .A(n254), .B(N8), .Y(n278) );
  AND2X2 U363 ( .A(n279), .B(n278), .Y(n338) );
  NAND2X1 U364 ( .A(n339), .B(n338), .Y(n286) );
  INVX2 U365 ( .A(\data[0][0] ), .Y(n282) );
  INVX2 U366 ( .A(w_data[0]), .Y(n370) );
  NAND3X1 U367 ( .A(n179), .B(n354), .C(n260), .Y(n281) );
  INVX2 U368 ( .A(n281), .Y(n287) );
  MUX2X1 U369 ( .B(n282), .A(n370), .S(n263), .Y(\nxt_data[0][0] ) );
  INVX2 U370 ( .A(\data[0][1] ), .Y(n283) );
  INVX2 U371 ( .A(w_data[1]), .Y(n372) );
  MUX2X1 U372 ( .B(n283), .A(n372), .S(n263), .Y(\nxt_data[0][1] ) );
  INVX2 U373 ( .A(\data[0][2] ), .Y(n284) );
  INVX2 U374 ( .A(w_data[2]), .Y(n374) );
  MUX2X1 U375 ( .B(n284), .A(n374), .S(n263), .Y(\nxt_data[0][2] ) );
  INVX2 U376 ( .A(\data[0][3] ), .Y(n285) );
  INVX2 U377 ( .A(w_data[3]), .Y(n376) );
  MUX2X1 U378 ( .B(n285), .A(n376), .S(n263), .Y(\nxt_data[0][3] ) );
  INVX2 U379 ( .A(\data[0][4] ), .Y(n288) );
  INVX2 U380 ( .A(w_data[4]), .Y(n378) );
  MUX2X1 U381 ( .B(n288), .A(n378), .S(n262), .Y(\nxt_data[0][4] ) );
  INVX2 U382 ( .A(\data[0][5] ), .Y(n289) );
  INVX2 U383 ( .A(w_data[5]), .Y(n380) );
  MUX2X1 U384 ( .B(n289), .A(n380), .S(n262), .Y(\nxt_data[0][5] ) );
  INVX2 U385 ( .A(\data[0][6] ), .Y(n290) );
  INVX2 U386 ( .A(w_data[6]), .Y(n382) );
  MUX2X1 U387 ( .B(n290), .A(n382), .S(n262), .Y(\nxt_data[0][6] ) );
  INVX2 U388 ( .A(\data[0][7] ), .Y(n291) );
  INVX2 U389 ( .A(w_data[7]), .Y(n384) );
  MUX2X1 U390 ( .B(n291), .A(n384), .S(n262), .Y(\nxt_data[0][7] ) );
  INVX2 U391 ( .A(\data[1][0] ), .Y(n293) );
  NAND3X1 U392 ( .A(n179), .B(n256), .C(n260), .Y(n292) );
  INVX2 U393 ( .A(n292), .Y(n297) );
  NAND2X1 U394 ( .A(n339), .B(n189), .Y(n307) );
  MUX2X1 U395 ( .B(n293), .A(n370), .S(n269), .Y(\nxt_data[1][0] ) );
  INVX2 U396 ( .A(\data[1][1] ), .Y(n294) );
  MUX2X1 U397 ( .B(n294), .A(n372), .S(n269), .Y(\nxt_data[1][1] ) );
  INVX2 U398 ( .A(\data[1][2] ), .Y(n295) );
  MUX2X1 U399 ( .B(n295), .A(n374), .S(n269), .Y(\nxt_data[1][2] ) );
  INVX2 U400 ( .A(\data[1][3] ), .Y(n296) );
  MUX2X1 U401 ( .B(n296), .A(n376), .S(n269), .Y(\nxt_data[1][3] ) );
  INVX2 U402 ( .A(\data[1][4] ), .Y(n298) );
  MUX2X1 U403 ( .B(n298), .A(n378), .S(n267), .Y(\nxt_data[1][4] ) );
  INVX2 U404 ( .A(\data[1][5] ), .Y(n299) );
  MUX2X1 U405 ( .B(n299), .A(n380), .S(n267), .Y(\nxt_data[1][5] ) );
  INVX2 U406 ( .A(\data[1][6] ), .Y(n300) );
  MUX2X1 U407 ( .B(n300), .A(n382), .S(n267), .Y(\nxt_data[1][6] ) );
  INVX2 U408 ( .A(\data[1][7] ), .Y(n301) );
  MUX2X1 U409 ( .B(n301), .A(n384), .S(n267), .Y(\nxt_data[1][7] ) );
  INVX2 U410 ( .A(\data[2][0] ), .Y(n303) );
  NAND3X1 U411 ( .A(n179), .B(n255), .C(n354), .Y(n302) );
  INVX2 U412 ( .A(n302), .Y(n308) );
  NAND2X1 U413 ( .A(n259), .B(n189), .Y(n317) );
  MUX2X1 U414 ( .B(n303), .A(n370), .S(n268), .Y(\nxt_data[2][0] ) );
  INVX2 U415 ( .A(\data[2][1] ), .Y(n304) );
  MUX2X1 U416 ( .B(n304), .A(n372), .S(n268), .Y(\nxt_data[2][1] ) );
  INVX2 U417 ( .A(\data[2][2] ), .Y(n305) );
  MUX2X1 U418 ( .B(n305), .A(n374), .S(n268), .Y(\nxt_data[2][2] ) );
  INVX2 U419 ( .A(\data[2][3] ), .Y(n306) );
  MUX2X1 U420 ( .B(n306), .A(n376), .S(n268), .Y(\nxt_data[2][3] ) );
  INVX2 U421 ( .A(\data[2][4] ), .Y(n309) );
  MUX2X1 U422 ( .B(n309), .A(n378), .S(n265), .Y(\nxt_data[2][4] ) );
  INVX2 U423 ( .A(\data[2][5] ), .Y(n310) );
  MUX2X1 U424 ( .B(n310), .A(n380), .S(n265), .Y(\nxt_data[2][5] ) );
  INVX2 U425 ( .A(\data[2][6] ), .Y(n311) );
  MUX2X1 U426 ( .B(n311), .A(n382), .S(n265), .Y(\nxt_data[2][6] ) );
  INVX2 U427 ( .A(\data[2][7] ), .Y(n312) );
  MUX2X1 U428 ( .B(n312), .A(n384), .S(n265), .Y(\nxt_data[2][7] ) );
  INVX2 U429 ( .A(\data[3][0] ), .Y(n313) );
  MUX2X1 U430 ( .B(n313), .A(n370), .S(n266), .Y(\nxt_data[3][0] ) );
  INVX2 U431 ( .A(\data[3][1] ), .Y(n314) );
  MUX2X1 U432 ( .B(n314), .A(n372), .S(n266), .Y(\nxt_data[3][1] ) );
  INVX2 U433 ( .A(\data[3][2] ), .Y(n315) );
  MUX2X1 U434 ( .B(n315), .A(n374), .S(n266), .Y(\nxt_data[3][2] ) );
  INVX2 U435 ( .A(\data[3][3] ), .Y(n316) );
  MUX2X1 U436 ( .B(n316), .A(n376), .S(n266), .Y(\nxt_data[3][3] ) );
  INVX2 U437 ( .A(\data[3][4] ), .Y(n318) );
  MUX2X1 U438 ( .B(n318), .A(n378), .S(n264), .Y(\nxt_data[3][4] ) );
  INVX2 U439 ( .A(\data[3][5] ), .Y(n319) );
  MUX2X1 U440 ( .B(n319), .A(n380), .S(n264), .Y(\nxt_data[3][5] ) );
  INVX2 U441 ( .A(\data[3][6] ), .Y(n320) );
  MUX2X1 U442 ( .B(n320), .A(n382), .S(n264), .Y(\nxt_data[3][6] ) );
  INVX2 U443 ( .A(\data[3][7] ), .Y(n321) );
  MUX2X1 U444 ( .B(n321), .A(n384), .S(n264), .Y(\nxt_data[3][7] ) );
  INVX2 U445 ( .A(\data[4][0] ), .Y(n324) );
  NAND3X1 U446 ( .A(n192), .B(n354), .C(n260), .Y(n322) );
  INVX2 U447 ( .A(n322), .Y(n329) );
  NAND2X1 U448 ( .A(n259), .B(n189), .Y(n346) );
  NAND2X1 U449 ( .A(n286), .B(n329), .Y(n323) );
  INVX2 U450 ( .A(n323), .Y(n327) );
  MUX2X1 U451 ( .B(n324), .A(n370), .S(n327), .Y(\nxt_data[4][0] ) );
  INVX2 U452 ( .A(\data[4][1] ), .Y(n325) );
  MUX2X1 U453 ( .B(n325), .A(n372), .S(n327), .Y(\nxt_data[4][1] ) );
  INVX2 U454 ( .A(\data[4][2] ), .Y(n326) );
  INVX2 U455 ( .A(\data[4][3] ), .Y(n328) );
  INVX2 U456 ( .A(\data[4][4] ), .Y(n331) );
  NAND2X1 U457 ( .A(n346), .B(n329), .Y(n330) );
  MUX2X1 U458 ( .B(n331), .A(n378), .S(n334), .Y(\nxt_data[4][4] ) );
  INVX2 U459 ( .A(\data[4][5] ), .Y(n332) );
  MUX2X1 U460 ( .B(n332), .A(n380), .S(n334), .Y(\nxt_data[4][5] ) );
  INVX2 U461 ( .A(\data[4][6] ), .Y(n333) );
  MUX2X1 U462 ( .B(n333), .A(n382), .S(n178), .Y(\nxt_data[4][6] ) );
  INVX2 U463 ( .A(\data[4][7] ), .Y(n335) );
  MUX2X1 U464 ( .B(n335), .A(n384), .S(n334), .Y(\nxt_data[4][7] ) );
  INVX2 U465 ( .A(\data[5][0] ), .Y(n341) );
  NAND3X1 U466 ( .A(n192), .B(n256), .C(n260), .Y(n337) );
  INVX2 U467 ( .A(n337), .Y(n347) );
  NAND2X1 U468 ( .A(n259), .B(n338), .Y(n361) );
  NAND2X1 U469 ( .A(n361), .B(n347), .Y(n340) );
  INVX2 U470 ( .A(n340), .Y(n344) );
  INVX2 U471 ( .A(\data[5][1] ), .Y(n342) );
  INVX2 U472 ( .A(\data[5][2] ), .Y(n343) );
  MUX2X1 U473 ( .B(n343), .A(n374), .S(n344), .Y(\nxt_data[5][2] ) );
  INVX2 U474 ( .A(\data[5][3] ), .Y(n345) );
  MUX2X1 U475 ( .B(n345), .A(n376), .S(n344), .Y(\nxt_data[5][3] ) );
  INVX2 U476 ( .A(\data[5][4] ), .Y(n349) );
  NAND2X1 U477 ( .A(n346), .B(n347), .Y(n348) );
  MUX2X1 U478 ( .B(n349), .A(n378), .S(n183), .Y(\nxt_data[5][4] ) );
  INVX2 U479 ( .A(\data[5][5] ), .Y(n350) );
  MUX2X1 U480 ( .B(n350), .A(n380), .S(n182), .Y(\nxt_data[5][5] ) );
  INVX2 U481 ( .A(\data[5][6] ), .Y(n351) );
  MUX2X1 U482 ( .B(n351), .A(n382), .S(n181), .Y(\nxt_data[5][6] ) );
  INVX2 U483 ( .A(\data[5][7] ), .Y(n353) );
  MUX2X1 U484 ( .B(n353), .A(n384), .S(n352), .Y(\nxt_data[5][7] ) );
  INVX2 U485 ( .A(\data[6][0] ), .Y(n357) );
  NAND3X1 U486 ( .A(n192), .B(n255), .C(n354), .Y(n355) );
  INVX2 U487 ( .A(n355), .Y(n362) );
  NAND2X1 U488 ( .A(n361), .B(n362), .Y(n356) );
  INVX2 U489 ( .A(\data[6][1] ), .Y(n358) );
  INVX2 U490 ( .A(\data[6][2] ), .Y(n359) );
  MUX2X1 U491 ( .B(n359), .A(n374), .S(n367), .Y(\nxt_data[6][2] ) );
  INVX2 U492 ( .A(\data[6][3] ), .Y(n360) );
  MUX2X1 U493 ( .B(n360), .A(n376), .S(n180), .Y(\nxt_data[6][3] ) );
  INVX2 U494 ( .A(\data[6][4] ), .Y(n364) );
  NAND2X1 U495 ( .A(n361), .B(n362), .Y(n363) );
  INVX2 U496 ( .A(n356), .Y(n367) );
  MUX2X1 U497 ( .B(n364), .A(n378), .S(n367), .Y(\nxt_data[6][4] ) );
  INVX2 U498 ( .A(\data[6][5] ), .Y(n365) );
  MUX2X1 U499 ( .B(n365), .A(n380), .S(n367), .Y(\nxt_data[6][5] ) );
  INVX2 U500 ( .A(\data[6][6] ), .Y(n366) );
  INVX2 U501 ( .A(\data[6][7] ), .Y(n368) );
  INVX2 U502 ( .A(\data[7][0] ), .Y(n371) );
  MUX2X1 U503 ( .B(n371), .A(n370), .S(n190), .Y(\nxt_data[7][0] ) );
  INVX2 U504 ( .A(\data[7][1] ), .Y(n373) );
  MUX2X1 U505 ( .B(n373), .A(n372), .S(n190), .Y(\nxt_data[7][1] ) );
  INVX2 U506 ( .A(\data[7][2] ), .Y(n375) );
  MUX2X1 U507 ( .B(n375), .A(n374), .S(n190), .Y(\nxt_data[7][2] ) );
  INVX2 U508 ( .A(\data[7][3] ), .Y(n377) );
  MUX2X1 U509 ( .B(n377), .A(n376), .S(n190), .Y(\nxt_data[7][3] ) );
  INVX2 U510 ( .A(\data[7][4] ), .Y(n379) );
  MUX2X1 U511 ( .B(n379), .A(n378), .S(n190), .Y(\nxt_data[7][4] ) );
  INVX2 U512 ( .A(\data[7][5] ), .Y(n381) );
  MUX2X1 U513 ( .B(n381), .A(n380), .S(n190), .Y(\nxt_data[7][5] ) );
  INVX2 U514 ( .A(\data[7][6] ), .Y(n383) );
  MUX2X1 U515 ( .B(n383), .A(n382), .S(n190), .Y(\nxt_data[7][6] ) );
  INVX2 U516 ( .A(\data[7][7] ), .Y(n385) );
  MUX2X1 U517 ( .B(n385), .A(n384), .S(n190), .Y(\nxt_data[7][7] ) );
endmodule

