// $Id: $
// File name:   upDownCounter.sv
// Created:     4/17/2015
// Author:      James Alliger
// Lab Section: 337-05
// Version:     1.0  Initial Design Entry
// Description: A counter that can count both up and down based on the inputs

module upDownCounter
#(
  parameter BITSIZE = 4 // the default is four bits. this is to make it easy to write
  )
( 
  input wire clk,
  input wire n_rst,
  input wire up,
  input wire down,
  output reg [BITSIZE - 1: 0]count_out
  
  );
  
  reg [BITSIZE - 1:0]nxt_count;
  
  always_ff @( posedge clk, negedge n_rst)
  begin
    if (n_rst ==1'b0)
      begin
        count_out <= '0;
      end
    else
      begin
        count_out <= nxt_count;
      end
    end
    
    always_comb
    begin
        nxt_count = count_out;
      if (up == down) //catch all for 1=1 and 0=0
        nxt_count = count_out;
      else if(up)
        nxt_count = count_out +1;
      else if(down & count_out)
        nxt_count = count_out -1;
    end
       
endmodule